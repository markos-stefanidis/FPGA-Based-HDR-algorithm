module g_green_lut(
	input clk,
	input clk_en,
	input [5:0] pixel,
	
	output reg [11:0] data
);

	always@(posedge clk) begin
		if(clk_en) begin
			case(pixel)
				6'h00: data <= 12'b000000000000;
				6'h01: data <= 12'b000000111011;
				6'h02: data <= 12'b000001110010;
				6'h03: data <= 12'b000010100101;
				6'h04: data <= 12'b000011010010;
				6'h05: data <= 12'b000011111100;
				6'h06: data <= 12'b000100100010;
				6'h07: data <= 12'b000101000010;
				6'h08: data <= 12'b000101011011;
				6'h09: data <= 12'b000101101111;
				6'h0A: data <= 12'b000110000000;
				6'h0B: data <= 12'b000110010001;
				6'h0C: data <= 12'b000110100001;
				6'h0D: data <= 12'b000110110010;
				6'h0E: data <= 12'b000111000011;
				6'h0F: data <= 12'b000111010101;
				6'h10: data <= 12'b000111100111;
				6'h11: data <= 12'b000111111001;
				6'h12: data <= 12'b001000001001;
				6'h13: data <= 12'b001000011001;
				6'h14: data <= 12'b001000101001;
				6'h15: data <= 12'b001000111000;
				6'h16: data <= 12'b001001000111;
				6'h17: data <= 12'b001001010101;
				6'h18: data <= 12'b001001100011;
				6'h19: data <= 12'b001001110001;
				6'h1A: data <= 12'b001001111110;
				6'h1B: data <= 12'b001010001010;
				6'h1C: data <= 12'b001010010111;
				6'h1D: data <= 12'b001010100011;
				6'h1E: data <= 12'b001010110000;
				6'h1F: data <= 12'b001010111101;
				6'h20: data <= 12'b001011001010;
				6'h21: data <= 12'b001011011000;
				6'h22: data <= 12'b001011100101;
				6'h23: data <= 12'b001011110010;
				6'h24: data <= 12'b001100000000;
				6'h25: data <= 12'b001100001110;
				6'h26: data <= 12'b001100011101;
				6'h27: data <= 12'b001100101100;
				6'h28: data <= 12'b001100111100;
				6'h29: data <= 12'b001101001100;
				6'h2A: data <= 12'b001101011100;
				6'h2B: data <= 12'b001101101100;
				6'h2C: data <= 12'b001101111100;
				6'h2D: data <= 12'b001110001010;
				6'h2E: data <= 12'b001110011001;
				6'h2F: data <= 12'b001110100111;
				6'h30: data <= 12'b001110110100;
				6'h31: data <= 12'b001111000001;
				6'h32: data <= 12'b001111001110;
				6'h33: data <= 12'b001111011010;
				6'h34: data <= 12'b001111100111;
				6'h35: data <= 12'b001111110011;
				6'h36: data <= 12'b001111111111;
				6'h37: data <= 12'b010000001011;
				6'h38: data <= 12'b010000011000;
				6'h39: data <= 12'b010000100101;
				6'h3A: data <= 12'b010000110001;
				6'h3B: data <= 12'b010000111100;
				6'h3C: data <= 12'b010001001000;
				6'h3D: data <= 12'b010001010011;
				6'h3E: data <= 12'b010001011110;
				6'h3F: data <= 12'b010001101000;
			endcase
		end
	end

endmodule
