module exp_lut(
	input clk,
	input clk_en,
	input [7:0] addr,

	output reg [31:0] data
);

	always@(posedge clk) begin
		if(clk_en) begin
			case(addr)
				8'd0:    data <= 32'b00000000000000000000000000010000;
				8'd1:    data <= 32'b00000000000000000000000000010001;
				8'd2:    data <= 32'b00000000000000000000000000010010;
				8'd3:    data <= 32'b00000000000000000000000000010011;
				8'd4:    data <= 32'b00000000000000000000000000010100;
				8'd5:    data <= 32'b00000000000000000000000000010101;
				8'd6:    data <= 32'b00000000000000000000000000010111;
				8'd7:    data <= 32'b00000000000000000000000000011000;
				8'd8:    data <= 32'b00000000000000000000000000011010;
				8'd9:    data <= 32'b00000000000000000000000000011100;
				8'd10:   data <= 32'b00000000000000000000000000011101;
				8'd11:   data <= 32'b00000000000000000000000000011111;
				8'd12:   data <= 32'b00000000000000000000000000100001;
				8'd13:   data <= 32'b00000000000000000000000000100100;
				8'd14:   data <= 32'b00000000000000000000000000100110;
				8'd15:   data <= 32'b00000000000000000000000000101000;
				8'd16:   data <= 32'b00000000000000000000000000101011;
				8'd17:   data <= 32'b00000000000000000000000000101110;
				8'd18:   data <= 32'b00000000000000000000000000110001;
				8'd19:   data <= 32'b00000000000000000000000000110100;
				8'd20:   data <= 32'b00000000000000000000000000110111;
				8'd21:   data <= 32'b00000000000000000000000000111011;
				8'd22:   data <= 32'b00000000000000000000000000111111;
				8'd23:   data <= 32'b00000000000000000000000001000011;
				8'd24:   data <= 32'b00000000000000000000000001000111;
				8'd25:   data <= 32'b00000000000000000000000001001100;
				8'd26:   data <= 32'b00000000000000000000000001010001;
				8'd27:   data <= 32'b00000000000000000000000001010110;
				8'd28:   data <= 32'b00000000000000000000000001011100;
				8'd29:   data <= 32'b00000000000000000000000001100010;
				8'd30:   data <= 32'b00000000000000000000000001101000;
				8'd31:   data <= 32'b00000000000000000000000001101111;
				8'd32:   data <= 32'b00000000000000000000000001110110;
				8'd33:   data <= 32'b00000000000000000000000001111101;
				8'd34:   data <= 32'b00000000000000000000000010000101;
				8'd35:   data <= 32'b00000000000000000000000010001110;
				8'd36:   data <= 32'b00000000000000000000000010010111;
				8'd37:   data <= 32'b00000000000000000000000010100001;
				8'd38:   data <= 32'b00000000000000000000000010101100;
				8'd39:   data <= 32'b00000000000000000000000010110111;
				8'd40:   data <= 32'b00000000000000000000000011000010;
				8'd41:   data <= 32'b00000000000000000000000011001111;
				8'd42:   data <= 32'b00000000000000000000000011011100;
				8'd43:   data <= 32'b00000000000000000000000011101011;
				8'd44:   data <= 32'b00000000000000000000000011111010;
				8'd45:   data <= 32'b00000000000000000000000100001010;
				8'd46:   data <= 32'b00000000000000000000000100011011;
				8'd47:   data <= 32'b00000000000000000000000100101101;
				8'd48:   data <= 32'b00000000000000000000000101000001;
				8'd49:   data <= 32'b00000000000000000000000101010110;
				8'd50:   data <= 32'b00000000000000000000000101101100;
				8'd51:   data <= 32'b00000000000000000000000110000011;
				8'd52:   data <= 32'b00000000000000000000000110011100;
				8'd53:   data <= 32'b00000000000000000000000110110111;
				8'd54:   data <= 32'b00000000000000000000000111010011;
				8'd55:   data <= 32'b00000000000000000000000111110001;
				8'd56:   data <= 32'b00000000000000000000001000010001;
				8'd57:   data <= 32'b00000000000000000000001000110100;
				8'd58:   data <= 32'b00000000000000000000001001011000;
				8'd59:   data <= 32'b00000000000000000000001001111111;
				8'd60:   data <= 32'b00000000000000000000001010101000;
				8'd61:   data <= 32'b00000000000000000000001011010100;
				8'd62:   data <= 32'b00000000000000000000001100000010;
				8'd63:   data <= 32'b00000000000000000000001100110100;
				8'd64:   data <= 32'b00000000000000000000001101101001;
				8'd65:   data <= 32'b00000000000000000000001110100001;
				8'd66:   data <= 32'b00000000000000000000001111011101;
				8'd67:   data <= 32'b00000000000000000000010000011101;
				8'd68:   data <= 32'b00000000000000000000010001100001;
				8'd69:   data <= 32'b00000000000000000000010010101010;
				8'd70:   data <= 32'b00000000000000000000010011110111;
				8'd71:   data <= 32'b00000000000000000000010101001001;
				8'd72:   data <= 32'b00000000000000000000010110100000;
				8'd73:   data <= 32'b00000000000000000000010111111101;
				8'd74:   data <= 32'b00000000000000000000011001100000;
				8'd75:   data <= 32'b00000000000000000000011011001001;
				8'd76:   data <= 32'b00000000000000000000011100111001;
				8'd77:   data <= 32'b00000000000000000000011110110000;
				8'd78:   data <= 32'b00000000000000000000100000101111;
				8'd79:   data <= 32'b00000000000000000000100010110110;
				8'd80:   data <= 32'b00000000000000000000100101000110;
				8'd81:   data <= 32'b00000000000000000000100111011111;
				8'd82:   data <= 32'b00000000000000000000101010000010;
				8'd83:   data <= 32'b00000000000000000000101100110000;
				8'd84:   data <= 32'b00000000000000000000101111101001;
				8'd85:   data <= 32'b00000000000000000000110010101101;
				8'd86:   data <= 32'b00000000000000000000110101111111;
				8'd87:   data <= 32'b00000000000000000000111001011101;
				8'd88:   data <= 32'b00000000000000000000111101001011;
				8'd89:   data <= 32'b00000000000000000001000001000111;
				8'd90:   data <= 32'b00000000000000000001000101010100;
				8'd91:   data <= 32'b00000000000000000001001001110010;
				8'd92:   data <= 32'b00000000000000000001001110100011;
				8'd93:   data <= 32'b00000000000000000001010011100111;
				8'd94:   data <= 32'b00000000000000000001011001000000;
				8'd95:   data <= 32'b00000000000000000001011110101111;
				8'd96:   data <= 32'b00000000000000000001100100110110;
				8'd97:   data <= 32'b00000000000000000001101011010111;
				8'd98:   data <= 32'b00000000000000000001110010010010;
				8'd99:   data <= 32'b00000000000000000001111001101010;
				8'd100:  data <= 32'b00000000000000000010000001100000;
				8'd101:  data <= 32'b00000000000000000010001001110110;
				8'd102:  data <= 32'b00000000000000000010010010101111;
				8'd103:  data <= 32'b00000000000000000010011100001101;
				8'd104:  data <= 32'b00000000000000000010100110010010;
				8'd105:  data <= 32'b00000000000000000010110001000000;
				8'd106:  data <= 32'b00000000000000000010111100011011;
				8'd107:  data <= 32'b00000000000000000011001000100101;
				8'd108:  data <= 32'b00000000000000000011010101100000;
				8'd109:  data <= 32'b00000000000000000011100011010010;
				8'd110:  data <= 32'b00000000000000000011110001111100;
				8'd111:  data <= 32'b00000000000000000100000001100011;
				8'd112:  data <= 32'b00000000000000000100010010001010;
				8'd113:  data <= 32'b00000000000000000100100011110101;
				8'd114:  data <= 32'b00000000000000000100110110101010;
				8'd115:  data <= 32'b00000000000000000101001010101100;
				8'd116:  data <= 32'b00000000000000000101100000000001;
				8'd117:  data <= 32'b00000000000000000101110110101110;
				8'd118:  data <= 32'b00000000000000000110001110111001;
				8'd119:  data <= 32'b00000000000000000110101000100111;
				8'd120:  data <= 32'b00000000000000000111000100000000;
				8'd121:  data <= 32'b00000000000000000111100001001010;
				8'd122:  data <= 32'b00000000000000001000000000001100;
				8'd123:  data <= 32'b00000000000000001000100001001110;
				8'd124:  data <= 32'b00000000000000001001000100011001;
				8'd125:  data <= 32'b00000000000000001001101001110100;
				8'd126:  data <= 32'b00000000000000001010010001101010;
				8'd127:  data <= 32'b00000000000000001010111100000101;
				8'd128:  data <= 32'b00000000000000001011101001001111;
				8'd129:  data <= 32'b00000000000000001100011001010011;
				8'd130:  data <= 32'b00000000000000001101001100011101;
				8'd131:  data <= 32'b00000000000000001110000010111011;
				8'd132:  data <= 32'b00000000000000001110111100111010;
				8'd133:  data <= 32'b00000000000000001111111010100111;
				8'd134:  data <= 32'b00000000000000010000111100010100;
				8'd135:  data <= 32'b00000000000000010010000010001111;
				8'd136:  data <= 32'b00000000000000010011001100101100;
				8'd137:  data <= 32'b00000000000000010100011011111011;
				8'd138:  data <= 32'b00000000000000010101110000010010;
				8'd139:  data <= 32'b00000000000000010111001010000101;
				8'd140:  data <= 32'b00000000000000011000101001101011;
				8'd141:  data <= 32'b00000000000000011010001111011011;
				8'd142:  data <= 32'b00000000000000011011111011101111;
				8'd143:  data <= 32'b00000000000000011101101111000010;
				8'd144:  data <= 32'b00000000000000011111101001110001;
				8'd145:  data <= 32'b00000000000000100001101100011011;
				8'd146:  data <= 32'b00000000000000100011110111011111;
				8'd147:  data <= 32'b00000000000000100110001011100010;
				8'd148:  data <= 32'b00000000000000101000101001001001;
				8'd149:  data <= 32'b00000000000000101011010000111001;
				8'd150:  data <= 32'b00000000000000101110000011011110;
				8'd151:  data <= 32'b00000000000000110001000001100100;
				8'd152:  data <= 32'b00000000000000110100001011111011;
				8'd153:  data <= 32'b00000000000000110111100011010101;
				8'd154:  data <= 32'b00000000000000111011001000101000;
				8'd155:  data <= 32'b00000000000000111110111100101110;
				8'd156:  data <= 32'b00000000000001000011000000100011;
				8'd157:  data <= 32'b00000000000001000111010101001001;
				8'd158:  data <= 32'b00000000000001001011111011100100;
				8'd159:  data <= 32'b00000000000001010000110100111111;
				8'd160:  data <= 32'b00000000000001010110000010100111;
				8'd161:  data <= 32'b00000000000001011011100101110000;
				8'd162:  data <= 32'b00000000000001100001011111110100;
				8'd163:  data <= 32'b00000000000001100111110010001111;
				8'd164:  data <= 32'b00000000000001101110011110101000;
				8'd165:  data <= 32'b00000000000001110101100110101001;
				8'd166:  data <= 32'b00000000000001111101001100000101;
				8'd167:  data <= 32'b00000000000010000101010000110100;
				8'd168:  data <= 32'b00000000000010001101110110111000;
				8'd169:  data <= 32'b00000000000010010111000000011010;
				8'd170:  data <= 32'b00000000000010100000101111101101;
				8'd171:  data <= 32'b00000000000010101011000111001101;
				8'd172:  data <= 32'b00000000000010110110001001100000;
				8'd173:  data <= 32'b00000000000011000001111001010110;
				8'd174:  data <= 32'b00000000000011001110011001101011;
				8'd175:  data <= 32'b00000000000011011011101101101000;
				8'd176:  data <= 32'b00000000000011101001111000100010;
				8'd177:  data <= 32'b00000000000011111000111101111011;
				8'd178:  data <= 32'b00000000000100001001000001100100;
				8'd179:  data <= 32'b00000000000100011010000111100000;
				8'd180:  data <= 32'b00000000000100101100010011111110;
				8'd181:  data <= 32'b00000000000100111111101011100011;
				8'd182:  data <= 32'b00000000000101010100010011000101;
				8'd183:  data <= 32'b00000000000101101010001111101110;
				8'd184:  data <= 32'b00000000000110000001100110111100;
				8'd185:  data <= 32'b00000000000110011010011110100110;
				8'd186:  data <= 32'b00000000000110110100111100111001;
				8'd187:  data <= 32'b00000000000111010001001000011111;
				8'd188:  data <= 32'b00000000000111101111001000011000;
				8'd189:  data <= 32'b00000000001000001111000100000111;
				8'd190:  data <= 32'b00000000001000110001000011101001;
				8'd191:  data <= 32'b00000000001001010101001111011111;
				8'd192:  data <= 32'b00000000001001111011110000101100;
				8'd193:  data <= 32'b00000000001010100100110000111001;
				8'd194:  data <= 32'b00000000001011010000011010010101;
				8'd195:  data <= 32'b00000000001011111110110111111100;
				8'd196:  data <= 32'b00000000001100110000010101010100;
				8'd197:  data <= 32'b00000000001101100100111110110110;
				8'd198:  data <= 32'b00000000001110011101000001101101;
				8'd199:  data <= 32'b00000000001111011000101011111000;
				8'd200:  data <= 32'b00000000010000011000001100010100;
				8'd201:  data <= 32'b00000000010001011011110010111000;
				8'd202:  data <= 32'b00000000010010100011110000011111;
				8'd203:  data <= 32'b00000000010011110000010111001000;
				8'd204:  data <= 32'b00000000010101000001111001111110;
				8'd205:  data <= 32'b00000000010110011000101101011001;
				8'd206:  data <= 32'b00000000010111110101000111000111;
				8'd207:  data <= 32'b00000000011001010111011110001110;
				8'd208:  data <= 32'b00000000011011000000001011010110;
				8'd209:  data <= 32'b00000000011100101111101000101001;
				8'd210:  data <= 32'b00000000011110100110010010000000;
				8'd211:  data <= 32'b00000000100000100100100101000110;
				8'd212:  data <= 32'b00000000100010101011000001100000;
				8'd213:  data <= 32'b00000000100100111010001000110110;
				8'd214:  data <= 32'b00000000100111010010011110111010;
				8'd215:  data <= 32'b00000000101001110100101001110100;
				8'd216:  data <= 32'b00000000101100100001010010000101;
				8'd217:  data <= 32'b00000000101111011001000010111010;
				8'd218:  data <= 32'b00000000110010011100101010010000;
				8'd219:  data <= 32'b00000000110101101100111001000001;
				8'd220:  data <= 32'b00000000111001001010100011010010;
				8'd221:  data <= 32'b00000000111100110110100000011111;
				8'd222:  data <= 32'b00000001000000110001101011101000;
				8'd223:  data <= 32'b00000001000100111101000011100010;
				8'd224:  data <= 32'b00000001001001011001101011000100;
				8'd225:  data <= 32'b00000001001110001000101001011001;
				8'd226:  data <= 32'b00000001010011001011001010010010;
				8'd227:  data <= 32'b00000001011000100010011110011010;
				8'd228:  data <= 32'b00000001011110001111111011100111;
				8'd229:  data <= 32'b00000001100100010100111101010010;
				8'd230:  data <= 32'b00000001101010110011000100101110;
				8'd231:  data <= 32'b00000001110001101011111001011111;
				8'd232:  data <= 32'b00000001111001000001001001110100;
				8'd233:  data <= 32'b00000010000000110100101011000011;
				8'd234:  data <= 32'b00000010001001001000011010001001;
				8'd235:  data <= 32'b00000010010001111110011100000011;
				8'd236:  data <= 32'b00000010011011011000111110010100;
				8'd237:  data <= 32'b00000010100101011010010111101001;
				8'd238:  data <= 32'b00000010110000000101001000011011;
				8'd239:  data <= 32'b00000010111011011011111011011001;
				8'd240:  data <= 32'b00000011000111100001100110010101;
				8'd241:  data <= 32'b00000011010100011001001010101110;
				8'd242:  data <= 32'b00000011100010000101110110011111;
				8'd243:  data <= 32'b00000011110000101011000100111010;
				8'd244:  data <= 32'b00000100000000001100011111010110;
				8'd245:  data <= 32'b00000100010000101101111110001111;
				8'd246:  data <= 32'b00000100100010010011101010000011;
				8'd247:  data <= 32'b00000100110101000001111100010010;
				8'd248:  data <= 32'b00000101001000111101100000100111;
				8'd249:  data <= 32'b00000101011110001011010110000010;
				8'd250:  data <= 32'b00000101110100110000110000000111;
				8'd251:  data <= 32'b00000110001100110011011000010101;
				8'd252:  data <= 32'b00000110100110011001001111011101;
				8'd253:  data <= 32'b00000111000001101000101111000101;
				8'd254:  data <= 32'b00000111011110101000101011010000;
				8'd255:  data <= 32'b00000111111101100000010100000100;
			endcase
		end
	end

endmodule
