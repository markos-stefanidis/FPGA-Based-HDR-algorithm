module exp_lut(
	input clk,
	input clk_en,
	input [11:0] address,
	
	output reg [31:0] data
);

	always@(posedge clk) begin
		if(clk_en) begin
			case(address)
				12'h000: data <= 32'b00000000000000000000000100000000;
				12'h001: data <= 32'b00000000000000000000000100000001;
				12'h002: data <= 32'b00000000000000000000000100000010;
				12'h003: data <= 32'b00000000000000000000000100000011;
				12'h004: data <= 32'b00000000000000000000000100000100;
				12'h005: data <= 32'b00000000000000000000000100000101;
				12'h006: data <= 32'b00000000000000000000000100000110;
				12'h007: data <= 32'b00000000000000000000000100000111;
				12'h008: data <= 32'b00000000000000000000000100001000;
				12'h009: data <= 32'b00000000000000000000000100001001;
				12'h00A: data <= 32'b00000000000000000000000100001010;
				12'h00B: data <= 32'b00000000000000000000000100001011;
				12'h00C: data <= 32'b00000000000000000000000100001100;
				12'h00D: data <= 32'b00000000000000000000000100001101;
				12'h00E: data <= 32'b00000000000000000000000100001110;
				12'h00F: data <= 32'b00000000000000000000000100001111;
				12'h010: data <= 32'b00000000000000000000000100010000;
				12'h011: data <= 32'b00000000000000000000000100010001;
				12'h012: data <= 32'b00000000000000000000000100010010;
				12'h013: data <= 32'b00000000000000000000000100010011;
				12'h014: data <= 32'b00000000000000000000000100010100;
				12'h015: data <= 32'b00000000000000000000000100010101;
				12'h016: data <= 32'b00000000000000000000000100010110;
				12'h017: data <= 32'b00000000000000000000000100011000;
				12'h018: data <= 32'b00000000000000000000000100011001;
				12'h019: data <= 32'b00000000000000000000000100011010;
				12'h01A: data <= 32'b00000000000000000000000100011011;
				12'h01B: data <= 32'b00000000000000000000000100011100;
				12'h01C: data <= 32'b00000000000000000000000100011101;
				12'h01D: data <= 32'b00000000000000000000000100011110;
				12'h01E: data <= 32'b00000000000000000000000100011111;
				12'h01F: data <= 32'b00000000000000000000000100100000;
				12'h020: data <= 32'b00000000000000000000000100100010;
				12'h021: data <= 32'b00000000000000000000000100100011;
				12'h022: data <= 32'b00000000000000000000000100100100;
				12'h023: data <= 32'b00000000000000000000000100100101;
				12'h024: data <= 32'b00000000000000000000000100100110;
				12'h025: data <= 32'b00000000000000000000000100100111;
				12'h026: data <= 32'b00000000000000000000000100101000;
				12'h027: data <= 32'b00000000000000000000000100101010;
				12'h028: data <= 32'b00000000000000000000000100101011;
				12'h029: data <= 32'b00000000000000000000000100101100;
				12'h02A: data <= 32'b00000000000000000000000100101101;
				12'h02B: data <= 32'b00000000000000000000000100101110;
				12'h02C: data <= 32'b00000000000000000000000100110000;
				12'h02D: data <= 32'b00000000000000000000000100110001;
				12'h02E: data <= 32'b00000000000000000000000100110010;
				12'h02F: data <= 32'b00000000000000000000000100110011;
				12'h030: data <= 32'b00000000000000000000000100110100;
				12'h031: data <= 32'b00000000000000000000000100110110;
				12'h032: data <= 32'b00000000000000000000000100110111;
				12'h033: data <= 32'b00000000000000000000000100111000;
				12'h034: data <= 32'b00000000000000000000000100111001;
				12'h035: data <= 32'b00000000000000000000000100111010;
				12'h036: data <= 32'b00000000000000000000000100111100;
				12'h037: data <= 32'b00000000000000000000000100111101;
				12'h038: data <= 32'b00000000000000000000000100111110;
				12'h039: data <= 32'b00000000000000000000000100111111;
				12'h03A: data <= 32'b00000000000000000000000101000001;
				12'h03B: data <= 32'b00000000000000000000000101000010;
				12'h03C: data <= 32'b00000000000000000000000101000011;
				12'h03D: data <= 32'b00000000000000000000000101000100;
				12'h03E: data <= 32'b00000000000000000000000101000110;
				12'h03F: data <= 32'b00000000000000000000000101000111;
				12'h040: data <= 32'b00000000000000000000000101001000;
				12'h041: data <= 32'b00000000000000000000000101001001;
				12'h042: data <= 32'b00000000000000000000000101001011;
				12'h043: data <= 32'b00000000000000000000000101001100;
				12'h044: data <= 32'b00000000000000000000000101001101;
				12'h045: data <= 32'b00000000000000000000000101001111;
				12'h046: data <= 32'b00000000000000000000000101010000;
				12'h047: data <= 32'b00000000000000000000000101010001;
				12'h048: data <= 32'b00000000000000000000000101010011;
				12'h049: data <= 32'b00000000000000000000000101010100;
				12'h04A: data <= 32'b00000000000000000000000101010101;
				12'h04B: data <= 32'b00000000000000000000000101010111;
				12'h04C: data <= 32'b00000000000000000000000101011000;
				12'h04D: data <= 32'b00000000000000000000000101011001;
				12'h04E: data <= 32'b00000000000000000000000101011011;
				12'h04F: data <= 32'b00000000000000000000000101011100;
				12'h050: data <= 32'b00000000000000000000000101011101;
				12'h051: data <= 32'b00000000000000000000000101011111;
				12'h052: data <= 32'b00000000000000000000000101100000;
				12'h053: data <= 32'b00000000000000000000000101100010;
				12'h054: data <= 32'b00000000000000000000000101100011;
				12'h055: data <= 32'b00000000000000000000000101100100;
				12'h056: data <= 32'b00000000000000000000000101100110;
				12'h057: data <= 32'b00000000000000000000000101100111;
				12'h058: data <= 32'b00000000000000000000000101101001;
				12'h059: data <= 32'b00000000000000000000000101101010;
				12'h05A: data <= 32'b00000000000000000000000101101011;
				12'h05B: data <= 32'b00000000000000000000000101101101;
				12'h05C: data <= 32'b00000000000000000000000101101110;
				12'h05D: data <= 32'b00000000000000000000000101110000;
				12'h05E: data <= 32'b00000000000000000000000101110001;
				12'h05F: data <= 32'b00000000000000000000000101110011;
				12'h060: data <= 32'b00000000000000000000000101110100;
				12'h061: data <= 32'b00000000000000000000000101110101;
				12'h062: data <= 32'b00000000000000000000000101110111;
				12'h063: data <= 32'b00000000000000000000000101111000;
				12'h064: data <= 32'b00000000000000000000000101111010;
				12'h065: data <= 32'b00000000000000000000000101111011;
				12'h066: data <= 32'b00000000000000000000000101111101;
				12'h067: data <= 32'b00000000000000000000000101111110;
				12'h068: data <= 32'b00000000000000000000000110000000;
				12'h069: data <= 32'b00000000000000000000000110000001;
				12'h06A: data <= 32'b00000000000000000000000110000011;
				12'h06B: data <= 32'b00000000000000000000000110000100;
				12'h06C: data <= 32'b00000000000000000000000110000110;
				12'h06D: data <= 32'b00000000000000000000000110000111;
				12'h06E: data <= 32'b00000000000000000000000110001001;
				12'h06F: data <= 32'b00000000000000000000000110001010;
				12'h070: data <= 32'b00000000000000000000000110001100;
				12'h071: data <= 32'b00000000000000000000000110001110;
				12'h072: data <= 32'b00000000000000000000000110001111;
				12'h073: data <= 32'b00000000000000000000000110010001;
				12'h074: data <= 32'b00000000000000000000000110010010;
				12'h075: data <= 32'b00000000000000000000000110010100;
				12'h076: data <= 32'b00000000000000000000000110010101;
				12'h077: data <= 32'b00000000000000000000000110010111;
				12'h078: data <= 32'b00000000000000000000000110011001;
				12'h079: data <= 32'b00000000000000000000000110011010;
				12'h07A: data <= 32'b00000000000000000000000110011100;
				12'h07B: data <= 32'b00000000000000000000000110011101;
				12'h07C: data <= 32'b00000000000000000000000110011111;
				12'h07D: data <= 32'b00000000000000000000000110100001;
				12'h07E: data <= 32'b00000000000000000000000110100010;
				12'h07F: data <= 32'b00000000000000000000000110100100;
				12'h080: data <= 32'b00000000000000000000000110100110;
				12'h081: data <= 32'b00000000000000000000000110100111;
				12'h082: data <= 32'b00000000000000000000000110101001;
				12'h083: data <= 32'b00000000000000000000000110101011;
				12'h084: data <= 32'b00000000000000000000000110101100;
				12'h085: data <= 32'b00000000000000000000000110101110;
				12'h086: data <= 32'b00000000000000000000000110110000;
				12'h087: data <= 32'b00000000000000000000000110110001;
				12'h088: data <= 32'b00000000000000000000000110110011;
				12'h089: data <= 32'b00000000000000000000000110110101;
				12'h08A: data <= 32'b00000000000000000000000110110110;
				12'h08B: data <= 32'b00000000000000000000000110111000;
				12'h08C: data <= 32'b00000000000000000000000110111010;
				12'h08D: data <= 32'b00000000000000000000000110111100;
				12'h08E: data <= 32'b00000000000000000000000110111101;
				12'h08F: data <= 32'b00000000000000000000000110111111;
				12'h090: data <= 32'b00000000000000000000000111000001;
				12'h091: data <= 32'b00000000000000000000000111000011;
				12'h092: data <= 32'b00000000000000000000000111000100;
				12'h093: data <= 32'b00000000000000000000000111000110;
				12'h094: data <= 32'b00000000000000000000000111001000;
				12'h095: data <= 32'b00000000000000000000000111001010;
				12'h096: data <= 32'b00000000000000000000000111001011;
				12'h097: data <= 32'b00000000000000000000000111001101;
				12'h098: data <= 32'b00000000000000000000000111001111;
				12'h099: data <= 32'b00000000000000000000000111010001;
				12'h09A: data <= 32'b00000000000000000000000111010011;
				12'h09B: data <= 32'b00000000000000000000000111010101;
				12'h09C: data <= 32'b00000000000000000000000111010110;
				12'h09D: data <= 32'b00000000000000000000000111011000;
				12'h09E: data <= 32'b00000000000000000000000111011010;
				12'h09F: data <= 32'b00000000000000000000000111011100;
				12'h0A0: data <= 32'b00000000000000000000000111011110;
				12'h0A1: data <= 32'b00000000000000000000000111100000;
				12'h0A2: data <= 32'b00000000000000000000000111100010;
				12'h0A3: data <= 32'b00000000000000000000000111100011;
				12'h0A4: data <= 32'b00000000000000000000000111100101;
				12'h0A5: data <= 32'b00000000000000000000000111100111;
				12'h0A6: data <= 32'b00000000000000000000000111101001;
				12'h0A7: data <= 32'b00000000000000000000000111101011;
				12'h0A8: data <= 32'b00000000000000000000000111101101;
				12'h0A9: data <= 32'b00000000000000000000000111101111;
				12'h0AA: data <= 32'b00000000000000000000000111110001;
				12'h0AB: data <= 32'b00000000000000000000000111110011;
				12'h0AC: data <= 32'b00000000000000000000000111110101;
				12'h0AD: data <= 32'b00000000000000000000000111110111;
				12'h0AE: data <= 32'b00000000000000000000000111111001;
				12'h0AF: data <= 32'b00000000000000000000000111111011;
				12'h0B0: data <= 32'b00000000000000000000000111111101;
				12'h0B1: data <= 32'b00000000000000000000000111111111;
				12'h0B2: data <= 32'b00000000000000000000001000000001;
				12'h0B3: data <= 32'b00000000000000000000001000000011;
				12'h0B4: data <= 32'b00000000000000000000001000000101;
				12'h0B5: data <= 32'b00000000000000000000001000000111;
				12'h0B6: data <= 32'b00000000000000000000001000001001;
				12'h0B7: data <= 32'b00000000000000000000001000001011;
				12'h0B8: data <= 32'b00000000000000000000001000001101;
				12'h0B9: data <= 32'b00000000000000000000001000001111;
				12'h0BA: data <= 32'b00000000000000000000001000010001;
				12'h0BB: data <= 32'b00000000000000000000001000010011;
				12'h0BC: data <= 32'b00000000000000000000001000010101;
				12'h0BD: data <= 32'b00000000000000000000001000010111;
				12'h0BE: data <= 32'b00000000000000000000001000011001;
				12'h0BF: data <= 32'b00000000000000000000001000011011;
				12'h0C0: data <= 32'b00000000000000000000001000011101;
				12'h0C1: data <= 32'b00000000000000000000001000100000;
				12'h0C2: data <= 32'b00000000000000000000001000100010;
				12'h0C3: data <= 32'b00000000000000000000001000100100;
				12'h0C4: data <= 32'b00000000000000000000001000100110;
				12'h0C5: data <= 32'b00000000000000000000001000101000;
				12'h0C6: data <= 32'b00000000000000000000001000101010;
				12'h0C7: data <= 32'b00000000000000000000001000101100;
				12'h0C8: data <= 32'b00000000000000000000001000101111;
				12'h0C9: data <= 32'b00000000000000000000001000110001;
				12'h0CA: data <= 32'b00000000000000000000001000110011;
				12'h0CB: data <= 32'b00000000000000000000001000110101;
				12'h0CC: data <= 32'b00000000000000000000001000110111;
				12'h0CD: data <= 32'b00000000000000000000001000111010;
				12'h0CE: data <= 32'b00000000000000000000001000111100;
				12'h0CF: data <= 32'b00000000000000000000001000111110;
				12'h0D0: data <= 32'b00000000000000000000001001000000;
				12'h0D1: data <= 32'b00000000000000000000001001000011;
				12'h0D2: data <= 32'b00000000000000000000001001000101;
				12'h0D3: data <= 32'b00000000000000000000001001000111;
				12'h0D4: data <= 32'b00000000000000000000001001001001;
				12'h0D5: data <= 32'b00000000000000000000001001001100;
				12'h0D6: data <= 32'b00000000000000000000001001001110;
				12'h0D7: data <= 32'b00000000000000000000001001010000;
				12'h0D8: data <= 32'b00000000000000000000001001010011;
				12'h0D9: data <= 32'b00000000000000000000001001010101;
				12'h0DA: data <= 32'b00000000000000000000001001010111;
				12'h0DB: data <= 32'b00000000000000000000001001011010;
				12'h0DC: data <= 32'b00000000000000000000001001011100;
				12'h0DD: data <= 32'b00000000000000000000001001011110;
				12'h0DE: data <= 32'b00000000000000000000001001100001;
				12'h0DF: data <= 32'b00000000000000000000001001100011;
				12'h0E0: data <= 32'b00000000000000000000001001100110;
				12'h0E1: data <= 32'b00000000000000000000001001101000;
				12'h0E2: data <= 32'b00000000000000000000001001101010;
				12'h0E3: data <= 32'b00000000000000000000001001101101;
				12'h0E4: data <= 32'b00000000000000000000001001101111;
				12'h0E5: data <= 32'b00000000000000000000001001110010;
				12'h0E6: data <= 32'b00000000000000000000001001110100;
				12'h0E7: data <= 32'b00000000000000000000001001110111;
				12'h0E8: data <= 32'b00000000000000000000001001111001;
				12'h0E9: data <= 32'b00000000000000000000001001111100;
				12'h0EA: data <= 32'b00000000000000000000001001111110;
				12'h0EB: data <= 32'b00000000000000000000001010000001;
				12'h0EC: data <= 32'b00000000000000000000001010000011;
				12'h0ED: data <= 32'b00000000000000000000001010000110;
				12'h0EE: data <= 32'b00000000000000000000001010001000;
				12'h0EF: data <= 32'b00000000000000000000001010001011;
				12'h0F0: data <= 32'b00000000000000000000001010001101;
				12'h0F1: data <= 32'b00000000000000000000001010010000;
				12'h0F2: data <= 32'b00000000000000000000001010010010;
				12'h0F3: data <= 32'b00000000000000000000001010010101;
				12'h0F4: data <= 32'b00000000000000000000001010011000;
				12'h0F5: data <= 32'b00000000000000000000001010011010;
				12'h0F6: data <= 32'b00000000000000000000001010011101;
				12'h0F7: data <= 32'b00000000000000000000001010011111;
				12'h0F8: data <= 32'b00000000000000000000001010100010;
				12'h0F9: data <= 32'b00000000000000000000001010100101;
				12'h0FA: data <= 32'b00000000000000000000001010100111;
				12'h0FB: data <= 32'b00000000000000000000001010101010;
				12'h0FC: data <= 32'b00000000000000000000001010101101;
				12'h0FD: data <= 32'b00000000000000000000001010101111;
				12'h0FE: data <= 32'b00000000000000000000001010110010;
				12'h0FF: data <= 32'b00000000000000000000001010110101;
				12'h100: data <= 32'b00000000000000000000001010110111;
				12'h101: data <= 32'b00000000000000000000001010111010;
				12'h102: data <= 32'b00000000000000000000001010111101;
				12'h103: data <= 32'b00000000000000000000001011000000;
				12'h104: data <= 32'b00000000000000000000001011000010;
				12'h105: data <= 32'b00000000000000000000001011000101;
				12'h106: data <= 32'b00000000000000000000001011001000;
				12'h107: data <= 32'b00000000000000000000001011001011;
				12'h108: data <= 32'b00000000000000000000001011001101;
				12'h109: data <= 32'b00000000000000000000001011010000;
				12'h10A: data <= 32'b00000000000000000000001011010011;
				12'h10B: data <= 32'b00000000000000000000001011010110;
				12'h10C: data <= 32'b00000000000000000000001011011001;
				12'h10D: data <= 32'b00000000000000000000001011011100;
				12'h10E: data <= 32'b00000000000000000000001011011110;
				12'h10F: data <= 32'b00000000000000000000001011100001;
				12'h110: data <= 32'b00000000000000000000001011100100;
				12'h111: data <= 32'b00000000000000000000001011100111;
				12'h112: data <= 32'b00000000000000000000001011101010;
				12'h113: data <= 32'b00000000000000000000001011101101;
				12'h114: data <= 32'b00000000000000000000001011110000;
				12'h115: data <= 32'b00000000000000000000001011110011;
				12'h116: data <= 32'b00000000000000000000001011110110;
				12'h117: data <= 32'b00000000000000000000001011111001;
				12'h118: data <= 32'b00000000000000000000001011111100;
				12'h119: data <= 32'b00000000000000000000001011111111;
				12'h11A: data <= 32'b00000000000000000000001100000010;
				12'h11B: data <= 32'b00000000000000000000001100000101;
				12'h11C: data <= 32'b00000000000000000000001100001000;
				12'h11D: data <= 32'b00000000000000000000001100001011;
				12'h11E: data <= 32'b00000000000000000000001100001110;
				12'h11F: data <= 32'b00000000000000000000001100010001;
				12'h120: data <= 32'b00000000000000000000001100010100;
				12'h121: data <= 32'b00000000000000000000001100010111;
				12'h122: data <= 32'b00000000000000000000001100011010;
				12'h123: data <= 32'b00000000000000000000001100011101;
				12'h124: data <= 32'b00000000000000000000001100100000;
				12'h125: data <= 32'b00000000000000000000001100100100;
				12'h126: data <= 32'b00000000000000000000001100100111;
				12'h127: data <= 32'b00000000000000000000001100101010;
				12'h128: data <= 32'b00000000000000000000001100101101;
				12'h129: data <= 32'b00000000000000000000001100110000;
				12'h12A: data <= 32'b00000000000000000000001100110011;
				12'h12B: data <= 32'b00000000000000000000001100110111;
				12'h12C: data <= 32'b00000000000000000000001100111010;
				12'h12D: data <= 32'b00000000000000000000001100111101;
				12'h12E: data <= 32'b00000000000000000000001101000000;
				12'h12F: data <= 32'b00000000000000000000001101000100;
				12'h130: data <= 32'b00000000000000000000001101000111;
				12'h131: data <= 32'b00000000000000000000001101001010;
				12'h132: data <= 32'b00000000000000000000001101001101;
				12'h133: data <= 32'b00000000000000000000001101010001;
				12'h134: data <= 32'b00000000000000000000001101010100;
				12'h135: data <= 32'b00000000000000000000001101010111;
				12'h136: data <= 32'b00000000000000000000001101011011;
				12'h137: data <= 32'b00000000000000000000001101011110;
				12'h138: data <= 32'b00000000000000000000001101100010;
				12'h139: data <= 32'b00000000000000000000001101100101;
				12'h13A: data <= 32'b00000000000000000000001101101000;
				12'h13B: data <= 32'b00000000000000000000001101101100;
				12'h13C: data <= 32'b00000000000000000000001101101111;
				12'h13D: data <= 32'b00000000000000000000001101110011;
				12'h13E: data <= 32'b00000000000000000000001101110110;
				12'h13F: data <= 32'b00000000000000000000001101111010;
				12'h140: data <= 32'b00000000000000000000001101111101;
				12'h141: data <= 32'b00000000000000000000001110000001;
				12'h142: data <= 32'b00000000000000000000001110000100;
				12'h143: data <= 32'b00000000000000000000001110001000;
				12'h144: data <= 32'b00000000000000000000001110001011;
				12'h145: data <= 32'b00000000000000000000001110001111;
				12'h146: data <= 32'b00000000000000000000001110010010;
				12'h147: data <= 32'b00000000000000000000001110010110;
				12'h148: data <= 32'b00000000000000000000001110011001;
				12'h149: data <= 32'b00000000000000000000001110011101;
				12'h14A: data <= 32'b00000000000000000000001110100001;
				12'h14B: data <= 32'b00000000000000000000001110100100;
				12'h14C: data <= 32'b00000000000000000000001110101000;
				12'h14D: data <= 32'b00000000000000000000001110101100;
				12'h14E: data <= 32'b00000000000000000000001110101111;
				12'h14F: data <= 32'b00000000000000000000001110110011;
				12'h150: data <= 32'b00000000000000000000001110110111;
				12'h151: data <= 32'b00000000000000000000001110111010;
				12'h152: data <= 32'b00000000000000000000001110111110;
				12'h153: data <= 32'b00000000000000000000001111000010;
				12'h154: data <= 32'b00000000000000000000001111000110;
				12'h155: data <= 32'b00000000000000000000001111001001;
				12'h156: data <= 32'b00000000000000000000001111001101;
				12'h157: data <= 32'b00000000000000000000001111010001;
				12'h158: data <= 32'b00000000000000000000001111010101;
				12'h159: data <= 32'b00000000000000000000001111011001;
				12'h15A: data <= 32'b00000000000000000000001111011101;
				12'h15B: data <= 32'b00000000000000000000001111100000;
				12'h15C: data <= 32'b00000000000000000000001111100100;
				12'h15D: data <= 32'b00000000000000000000001111101000;
				12'h15E: data <= 32'b00000000000000000000001111101100;
				12'h15F: data <= 32'b00000000000000000000001111110000;
				12'h160: data <= 32'b00000000000000000000001111110100;
				12'h161: data <= 32'b00000000000000000000001111111000;
				12'h162: data <= 32'b00000000000000000000001111111100;
				12'h163: data <= 32'b00000000000000000000010000000000;
				12'h164: data <= 32'b00000000000000000000010000000100;
				12'h165: data <= 32'b00000000000000000000010000001000;
				12'h166: data <= 32'b00000000000000000000010000001100;
				12'h167: data <= 32'b00000000000000000000010000010000;
				12'h168: data <= 32'b00000000000000000000010000010100;
				12'h169: data <= 32'b00000000000000000000010000011000;
				12'h16A: data <= 32'b00000000000000000000010000011100;
				12'h16B: data <= 32'b00000000000000000000010000100000;
				12'h16C: data <= 32'b00000000000000000000010000100101;
				12'h16D: data <= 32'b00000000000000000000010000101001;
				12'h16E: data <= 32'b00000000000000000000010000101101;
				12'h16F: data <= 32'b00000000000000000000010000110001;
				12'h170: data <= 32'b00000000000000000000010000110101;
				12'h171: data <= 32'b00000000000000000000010000111010;
				12'h172: data <= 32'b00000000000000000000010000111110;
				12'h173: data <= 32'b00000000000000000000010001000010;
				12'h174: data <= 32'b00000000000000000000010001000110;
				12'h175: data <= 32'b00000000000000000000010001001011;
				12'h176: data <= 32'b00000000000000000000010001001111;
				12'h177: data <= 32'b00000000000000000000010001010011;
				12'h178: data <= 32'b00000000000000000000010001011000;
				12'h179: data <= 32'b00000000000000000000010001011100;
				12'h17A: data <= 32'b00000000000000000000010001100000;
				12'h17B: data <= 32'b00000000000000000000010001100101;
				12'h17C: data <= 32'b00000000000000000000010001101001;
				12'h17D: data <= 32'b00000000000000000000010001101101;
				12'h17E: data <= 32'b00000000000000000000010001110010;
				12'h17F: data <= 32'b00000000000000000000010001110110;
				12'h180: data <= 32'b00000000000000000000010001111011;
				12'h181: data <= 32'b00000000000000000000010001111111;
				12'h182: data <= 32'b00000000000000000000010010000100;
				12'h183: data <= 32'b00000000000000000000010010001000;
				12'h184: data <= 32'b00000000000000000000010010001101;
				12'h185: data <= 32'b00000000000000000000010010010001;
				12'h186: data <= 32'b00000000000000000000010010010110;
				12'h187: data <= 32'b00000000000000000000010010011011;
				12'h188: data <= 32'b00000000000000000000010010011111;
				12'h189: data <= 32'b00000000000000000000010010100100;
				12'h18A: data <= 32'b00000000000000000000010010101001;
				12'h18B: data <= 32'b00000000000000000000010010101101;
				12'h18C: data <= 32'b00000000000000000000010010110010;
				12'h18D: data <= 32'b00000000000000000000010010110111;
				12'h18E: data <= 32'b00000000000000000000010010111011;
				12'h18F: data <= 32'b00000000000000000000010011000000;
				12'h190: data <= 32'b00000000000000000000010011000101;
				12'h191: data <= 32'b00000000000000000000010011001010;
				12'h192: data <= 32'b00000000000000000000010011001110;
				12'h193: data <= 32'b00000000000000000000010011010011;
				12'h194: data <= 32'b00000000000000000000010011011000;
				12'h195: data <= 32'b00000000000000000000010011011101;
				12'h196: data <= 32'b00000000000000000000010011100010;
				12'h197: data <= 32'b00000000000000000000010011100111;
				12'h198: data <= 32'b00000000000000000000010011101100;
				12'h199: data <= 32'b00000000000000000000010011110001;
				12'h19A: data <= 32'b00000000000000000000010011110101;
				12'h19B: data <= 32'b00000000000000000000010011111010;
				12'h19C: data <= 32'b00000000000000000000010011111111;
				12'h19D: data <= 32'b00000000000000000000010100000100;
				12'h19E: data <= 32'b00000000000000000000010100001001;
				12'h19F: data <= 32'b00000000000000000000010100001111;
				12'h1A0: data <= 32'b00000000000000000000010100010100;
				12'h1A1: data <= 32'b00000000000000000000010100011001;
				12'h1A2: data <= 32'b00000000000000000000010100011110;
				12'h1A3: data <= 32'b00000000000000000000010100100011;
				12'h1A4: data <= 32'b00000000000000000000010100101000;
				12'h1A5: data <= 32'b00000000000000000000010100101101;
				12'h1A6: data <= 32'b00000000000000000000010100110010;
				12'h1A7: data <= 32'b00000000000000000000010100111000;
				12'h1A8: data <= 32'b00000000000000000000010100111101;
				12'h1A9: data <= 32'b00000000000000000000010101000010;
				12'h1AA: data <= 32'b00000000000000000000010101000111;
				12'h1AB: data <= 32'b00000000000000000000010101001101;
				12'h1AC: data <= 32'b00000000000000000000010101010010;
				12'h1AD: data <= 32'b00000000000000000000010101010111;
				12'h1AE: data <= 32'b00000000000000000000010101011101;
				12'h1AF: data <= 32'b00000000000000000000010101100010;
				12'h1B0: data <= 32'b00000000000000000000010101100111;
				12'h1B1: data <= 32'b00000000000000000000010101101101;
				12'h1B2: data <= 32'b00000000000000000000010101110010;
				12'h1B3: data <= 32'b00000000000000000000010101111000;
				12'h1B4: data <= 32'b00000000000000000000010101111101;
				12'h1B5: data <= 32'b00000000000000000000010110000011;
				12'h1B6: data <= 32'b00000000000000000000010110001000;
				12'h1B7: data <= 32'b00000000000000000000010110001110;
				12'h1B8: data <= 32'b00000000000000000000010110010011;
				12'h1B9: data <= 32'b00000000000000000000010110011001;
				12'h1BA: data <= 32'b00000000000000000000010110011111;
				12'h1BB: data <= 32'b00000000000000000000010110100100;
				12'h1BC: data <= 32'b00000000000000000000010110101010;
				12'h1BD: data <= 32'b00000000000000000000010110110000;
				12'h1BE: data <= 32'b00000000000000000000010110110101;
				12'h1BF: data <= 32'b00000000000000000000010110111011;
				12'h1C0: data <= 32'b00000000000000000000010111000001;
				12'h1C1: data <= 32'b00000000000000000000010111000110;
				12'h1C2: data <= 32'b00000000000000000000010111001100;
				12'h1C3: data <= 32'b00000000000000000000010111010010;
				12'h1C4: data <= 32'b00000000000000000000010111011000;
				12'h1C5: data <= 32'b00000000000000000000010111011110;
				12'h1C6: data <= 32'b00000000000000000000010111100100;
				12'h1C7: data <= 32'b00000000000000000000010111101010;
				12'h1C8: data <= 32'b00000000000000000000010111101111;
				12'h1C9: data <= 32'b00000000000000000000010111110101;
				12'h1CA: data <= 32'b00000000000000000000010111111011;
				12'h1CB: data <= 32'b00000000000000000000011000000001;
				12'h1CC: data <= 32'b00000000000000000000011000000111;
				12'h1CD: data <= 32'b00000000000000000000011000001101;
				12'h1CE: data <= 32'b00000000000000000000011000010011;
				12'h1CF: data <= 32'b00000000000000000000011000011010;
				12'h1D0: data <= 32'b00000000000000000000011000100000;
				12'h1D1: data <= 32'b00000000000000000000011000100110;
				12'h1D2: data <= 32'b00000000000000000000011000101100;
				12'h1D3: data <= 32'b00000000000000000000011000110010;
				12'h1D4: data <= 32'b00000000000000000000011000111000;
				12'h1D5: data <= 32'b00000000000000000000011000111111;
				12'h1D6: data <= 32'b00000000000000000000011001000101;
				12'h1D7: data <= 32'b00000000000000000000011001001011;
				12'h1D8: data <= 32'b00000000000000000000011001010001;
				12'h1D9: data <= 32'b00000000000000000000011001011000;
				12'h1DA: data <= 32'b00000000000000000000011001011110;
				12'h1DB: data <= 32'b00000000000000000000011001100101;
				12'h1DC: data <= 32'b00000000000000000000011001101011;
				12'h1DD: data <= 32'b00000000000000000000011001110001;
				12'h1DE: data <= 32'b00000000000000000000011001111000;
				12'h1DF: data <= 32'b00000000000000000000011001111110;
				12'h1E0: data <= 32'b00000000000000000000011010000101;
				12'h1E1: data <= 32'b00000000000000000000011010001011;
				12'h1E2: data <= 32'b00000000000000000000011010010010;
				12'h1E3: data <= 32'b00000000000000000000011010011001;
				12'h1E4: data <= 32'b00000000000000000000011010011111;
				12'h1E5: data <= 32'b00000000000000000000011010100110;
				12'h1E6: data <= 32'b00000000000000000000011010101100;
				12'h1E7: data <= 32'b00000000000000000000011010110011;
				12'h1E8: data <= 32'b00000000000000000000011010111010;
				12'h1E9: data <= 32'b00000000000000000000011011000001;
				12'h1EA: data <= 32'b00000000000000000000011011000111;
				12'h1EB: data <= 32'b00000000000000000000011011001110;
				12'h1EC: data <= 32'b00000000000000000000011011010101;
				12'h1ED: data <= 32'b00000000000000000000011011011100;
				12'h1EE: data <= 32'b00000000000000000000011011100011;
				12'h1EF: data <= 32'b00000000000000000000011011101010;
				12'h1F0: data <= 32'b00000000000000000000011011110000;
				12'h1F1: data <= 32'b00000000000000000000011011110111;
				12'h1F2: data <= 32'b00000000000000000000011011111110;
				12'h1F3: data <= 32'b00000000000000000000011100000101;
				12'h1F4: data <= 32'b00000000000000000000011100001100;
				12'h1F5: data <= 32'b00000000000000000000011100010100;
				12'h1F6: data <= 32'b00000000000000000000011100011011;
				12'h1F7: data <= 32'b00000000000000000000011100100010;
				12'h1F8: data <= 32'b00000000000000000000011100101001;
				12'h1F9: data <= 32'b00000000000000000000011100110000;
				12'h1FA: data <= 32'b00000000000000000000011100110111;
				12'h1FB: data <= 32'b00000000000000000000011100111111;
				12'h1FC: data <= 32'b00000000000000000000011101000110;
				12'h1FD: data <= 32'b00000000000000000000011101001101;
				12'h1FE: data <= 32'b00000000000000000000011101010100;
				12'h1FF: data <= 32'b00000000000000000000011101011100;
				12'h200: data <= 32'b00000000000000000000011101100011;
				12'h201: data <= 32'b00000000000000000000011101101011;
				12'h202: data <= 32'b00000000000000000000011101110010;
				12'h203: data <= 32'b00000000000000000000011101111001;
				12'h204: data <= 32'b00000000000000000000011110000001;
				12'h205: data <= 32'b00000000000000000000011110001000;
				12'h206: data <= 32'b00000000000000000000011110010000;
				12'h207: data <= 32'b00000000000000000000011110011000;
				12'h208: data <= 32'b00000000000000000000011110011111;
				12'h209: data <= 32'b00000000000000000000011110100111;
				12'h20A: data <= 32'b00000000000000000000011110101110;
				12'h20B: data <= 32'b00000000000000000000011110110110;
				12'h20C: data <= 32'b00000000000000000000011110111110;
				12'h20D: data <= 32'b00000000000000000000011111000110;
				12'h20E: data <= 32'b00000000000000000000011111001101;
				12'h20F: data <= 32'b00000000000000000000011111010101;
				12'h210: data <= 32'b00000000000000000000011111011101;
				12'h211: data <= 32'b00000000000000000000011111100101;
				12'h212: data <= 32'b00000000000000000000011111101101;
				12'h213: data <= 32'b00000000000000000000011111110101;
				12'h214: data <= 32'b00000000000000000000011111111101;
				12'h215: data <= 32'b00000000000000000000100000000101;
				12'h216: data <= 32'b00000000000000000000100000001101;
				12'h217: data <= 32'b00000000000000000000100000010101;
				12'h218: data <= 32'b00000000000000000000100000011101;
				12'h219: data <= 32'b00000000000000000000100000100101;
				12'h21A: data <= 32'b00000000000000000000100000101101;
				12'h21B: data <= 32'b00000000000000000000100000110110;
				12'h21C: data <= 32'b00000000000000000000100000111110;
				12'h21D: data <= 32'b00000000000000000000100001000110;
				12'h21E: data <= 32'b00000000000000000000100001001110;
				12'h21F: data <= 32'b00000000000000000000100001010111;
				12'h220: data <= 32'b00000000000000000000100001011111;
				12'h221: data <= 32'b00000000000000000000100001100111;
				12'h222: data <= 32'b00000000000000000000100001110000;
				12'h223: data <= 32'b00000000000000000000100001111000;
				12'h224: data <= 32'b00000000000000000000100010000001;
				12'h225: data <= 32'b00000000000000000000100010001001;
				12'h226: data <= 32'b00000000000000000000100010010010;
				12'h227: data <= 32'b00000000000000000000100010011010;
				12'h228: data <= 32'b00000000000000000000100010100011;
				12'h229: data <= 32'b00000000000000000000100010101100;
				12'h22A: data <= 32'b00000000000000000000100010110100;
				12'h22B: data <= 32'b00000000000000000000100010111101;
				12'h22C: data <= 32'b00000000000000000000100011000110;
				12'h22D: data <= 32'b00000000000000000000100011001111;
				12'h22E: data <= 32'b00000000000000000000100011010111;
				12'h22F: data <= 32'b00000000000000000000100011100000;
				12'h230: data <= 32'b00000000000000000000100011101001;
				12'h231: data <= 32'b00000000000000000000100011110010;
				12'h232: data <= 32'b00000000000000000000100011111011;
				12'h233: data <= 32'b00000000000000000000100100000100;
				12'h234: data <= 32'b00000000000000000000100100001101;
				12'h235: data <= 32'b00000000000000000000100100010110;
				12'h236: data <= 32'b00000000000000000000100100011111;
				12'h237: data <= 32'b00000000000000000000100100101000;
				12'h238: data <= 32'b00000000000000000000100100110010;
				12'h239: data <= 32'b00000000000000000000100100111011;
				12'h23A: data <= 32'b00000000000000000000100101000100;
				12'h23B: data <= 32'b00000000000000000000100101001101;
				12'h23C: data <= 32'b00000000000000000000100101010111;
				12'h23D: data <= 32'b00000000000000000000100101100000;
				12'h23E: data <= 32'b00000000000000000000100101101001;
				12'h23F: data <= 32'b00000000000000000000100101110011;
				12'h240: data <= 32'b00000000000000000000100101111100;
				12'h241: data <= 32'b00000000000000000000100110000110;
				12'h242: data <= 32'b00000000000000000000100110001111;
				12'h243: data <= 32'b00000000000000000000100110011001;
				12'h244: data <= 32'b00000000000000000000100110100011;
				12'h245: data <= 32'b00000000000000000000100110101100;
				12'h246: data <= 32'b00000000000000000000100110110110;
				12'h247: data <= 32'b00000000000000000000100111000000;
				12'h248: data <= 32'b00000000000000000000100111001001;
				12'h249: data <= 32'b00000000000000000000100111010011;
				12'h24A: data <= 32'b00000000000000000000100111011101;
				12'h24B: data <= 32'b00000000000000000000100111100111;
				12'h24C: data <= 32'b00000000000000000000100111110001;
				12'h24D: data <= 32'b00000000000000000000100111111011;
				12'h24E: data <= 32'b00000000000000000000101000000101;
				12'h24F: data <= 32'b00000000000000000000101000001111;
				12'h250: data <= 32'b00000000000000000000101000011001;
				12'h251: data <= 32'b00000000000000000000101000100011;
				12'h252: data <= 32'b00000000000000000000101000101101;
				12'h253: data <= 32'b00000000000000000000101000110111;
				12'h254: data <= 32'b00000000000000000000101001000010;
				12'h255: data <= 32'b00000000000000000000101001001100;
				12'h256: data <= 32'b00000000000000000000101001010110;
				12'h257: data <= 32'b00000000000000000000101001100001;
				12'h258: data <= 32'b00000000000000000000101001101011;
				12'h259: data <= 32'b00000000000000000000101001110110;
				12'h25A: data <= 32'b00000000000000000000101010000000;
				12'h25B: data <= 32'b00000000000000000000101010001011;
				12'h25C: data <= 32'b00000000000000000000101010010101;
				12'h25D: data <= 32'b00000000000000000000101010100000;
				12'h25E: data <= 32'b00000000000000000000101010101010;
				12'h25F: data <= 32'b00000000000000000000101010110101;
				12'h260: data <= 32'b00000000000000000000101011000000;
				12'h261: data <= 32'b00000000000000000000101011001011;
				12'h262: data <= 32'b00000000000000000000101011010101;
				12'h263: data <= 32'b00000000000000000000101011100000;
				12'h264: data <= 32'b00000000000000000000101011101011;
				12'h265: data <= 32'b00000000000000000000101011110110;
				12'h266: data <= 32'b00000000000000000000101100000001;
				12'h267: data <= 32'b00000000000000000000101100001100;
				12'h268: data <= 32'b00000000000000000000101100010111;
				12'h269: data <= 32'b00000000000000000000101100100010;
				12'h26A: data <= 32'b00000000000000000000101100101101;
				12'h26B: data <= 32'b00000000000000000000101100111001;
				12'h26C: data <= 32'b00000000000000000000101101000100;
				12'h26D: data <= 32'b00000000000000000000101101001111;
				12'h26E: data <= 32'b00000000000000000000101101011010;
				12'h26F: data <= 32'b00000000000000000000101101100110;
				12'h270: data <= 32'b00000000000000000000101101110001;
				12'h271: data <= 32'b00000000000000000000101101111101;
				12'h272: data <= 32'b00000000000000000000101110001000;
				12'h273: data <= 32'b00000000000000000000101110010100;
				12'h274: data <= 32'b00000000000000000000101110011111;
				12'h275: data <= 32'b00000000000000000000101110101011;
				12'h276: data <= 32'b00000000000000000000101110110111;
				12'h277: data <= 32'b00000000000000000000101111000010;
				12'h278: data <= 32'b00000000000000000000101111001110;
				12'h279: data <= 32'b00000000000000000000101111011010;
				12'h27A: data <= 32'b00000000000000000000101111100110;
				12'h27B: data <= 32'b00000000000000000000101111110010;
				12'h27C: data <= 32'b00000000000000000000101111111110;
				12'h27D: data <= 32'b00000000000000000000110000001010;
				12'h27E: data <= 32'b00000000000000000000110000010110;
				12'h27F: data <= 32'b00000000000000000000110000100010;
				12'h280: data <= 32'b00000000000000000000110000101110;
				12'h281: data <= 32'b00000000000000000000110000111010;
				12'h282: data <= 32'b00000000000000000000110001000111;
				12'h283: data <= 32'b00000000000000000000110001010011;
				12'h284: data <= 32'b00000000000000000000110001011111;
				12'h285: data <= 32'b00000000000000000000110001101100;
				12'h286: data <= 32'b00000000000000000000110001111000;
				12'h287: data <= 32'b00000000000000000000110010000101;
				12'h288: data <= 32'b00000000000000000000110010010001;
				12'h289: data <= 32'b00000000000000000000110010011110;
				12'h28A: data <= 32'b00000000000000000000110010101010;
				12'h28B: data <= 32'b00000000000000000000110010110111;
				12'h28C: data <= 32'b00000000000000000000110011000100;
				12'h28D: data <= 32'b00000000000000000000110011010001;
				12'h28E: data <= 32'b00000000000000000000110011011110;
				12'h28F: data <= 32'b00000000000000000000110011101010;
				12'h290: data <= 32'b00000000000000000000110011110111;
				12'h291: data <= 32'b00000000000000000000110100000100;
				12'h292: data <= 32'b00000000000000000000110100010001;
				12'h293: data <= 32'b00000000000000000000110100011110;
				12'h294: data <= 32'b00000000000000000000110100101100;
				12'h295: data <= 32'b00000000000000000000110100111001;
				12'h296: data <= 32'b00000000000000000000110101000110;
				12'h297: data <= 32'b00000000000000000000110101010011;
				12'h298: data <= 32'b00000000000000000000110101100001;
				12'h299: data <= 32'b00000000000000000000110101101110;
				12'h29A: data <= 32'b00000000000000000000110101111100;
				12'h29B: data <= 32'b00000000000000000000110110001001;
				12'h29C: data <= 32'b00000000000000000000110110010111;
				12'h29D: data <= 32'b00000000000000000000110110100100;
				12'h29E: data <= 32'b00000000000000000000110110110010;
				12'h29F: data <= 32'b00000000000000000000110111000000;
				12'h2A0: data <= 32'b00000000000000000000110111001101;
				12'h2A1: data <= 32'b00000000000000000000110111011011;
				12'h2A2: data <= 32'b00000000000000000000110111101001;
				12'h2A3: data <= 32'b00000000000000000000110111110111;
				12'h2A4: data <= 32'b00000000000000000000111000000101;
				12'h2A5: data <= 32'b00000000000000000000111000010011;
				12'h2A6: data <= 32'b00000000000000000000111000100001;
				12'h2A7: data <= 32'b00000000000000000000111000101111;
				12'h2A8: data <= 32'b00000000000000000000111000111110;
				12'h2A9: data <= 32'b00000000000000000000111001001100;
				12'h2AA: data <= 32'b00000000000000000000111001011010;
				12'h2AB: data <= 32'b00000000000000000000111001101001;
				12'h2AC: data <= 32'b00000000000000000000111001110111;
				12'h2AD: data <= 32'b00000000000000000000111010000110;
				12'h2AE: data <= 32'b00000000000000000000111010010100;
				12'h2AF: data <= 32'b00000000000000000000111010100011;
				12'h2B0: data <= 32'b00000000000000000000111010110001;
				12'h2B1: data <= 32'b00000000000000000000111011000000;
				12'h2B2: data <= 32'b00000000000000000000111011001111;
				12'h2B3: data <= 32'b00000000000000000000111011011110;
				12'h2B4: data <= 32'b00000000000000000000111011101101;
				12'h2B5: data <= 32'b00000000000000000000111011111100;
				12'h2B6: data <= 32'b00000000000000000000111100001011;
				12'h2B7: data <= 32'b00000000000000000000111100011010;
				12'h2B8: data <= 32'b00000000000000000000111100101001;
				12'h2B9: data <= 32'b00000000000000000000111100111000;
				12'h2BA: data <= 32'b00000000000000000000111101000111;
				12'h2BB: data <= 32'b00000000000000000000111101010111;
				12'h2BC: data <= 32'b00000000000000000000111101100110;
				12'h2BD: data <= 32'b00000000000000000000111101110101;
				12'h2BE: data <= 32'b00000000000000000000111110000101;
				12'h2BF: data <= 32'b00000000000000000000111110010100;
				12'h2C0: data <= 32'b00000000000000000000111110100100;
				12'h2C1: data <= 32'b00000000000000000000111110110100;
				12'h2C2: data <= 32'b00000000000000000000111111000011;
				12'h2C3: data <= 32'b00000000000000000000111111010011;
				12'h2C4: data <= 32'b00000000000000000000111111100011;
				12'h2C5: data <= 32'b00000000000000000000111111110011;
				12'h2C6: data <= 32'b00000000000000000001000000000011;
				12'h2C7: data <= 32'b00000000000000000001000000010011;
				12'h2C8: data <= 32'b00000000000000000001000000100011;
				12'h2C9: data <= 32'b00000000000000000001000000110011;
				12'h2CA: data <= 32'b00000000000000000001000001000100;
				12'h2CB: data <= 32'b00000000000000000001000001010100;
				12'h2CC: data <= 32'b00000000000000000001000001100100;
				12'h2CD: data <= 32'b00000000000000000001000001110101;
				12'h2CE: data <= 32'b00000000000000000001000010000101;
				12'h2CF: data <= 32'b00000000000000000001000010010110;
				12'h2D0: data <= 32'b00000000000000000001000010100110;
				12'h2D1: data <= 32'b00000000000000000001000010110111;
				12'h2D2: data <= 32'b00000000000000000001000011001000;
				12'h2D3: data <= 32'b00000000000000000001000011011001;
				12'h2D4: data <= 32'b00000000000000000001000011101001;
				12'h2D5: data <= 32'b00000000000000000001000011111010;
				12'h2D6: data <= 32'b00000000000000000001000100001011;
				12'h2D7: data <= 32'b00000000000000000001000100011100;
				12'h2D8: data <= 32'b00000000000000000001000100101110;
				12'h2D9: data <= 32'b00000000000000000001000100111111;
				12'h2DA: data <= 32'b00000000000000000001000101010000;
				12'h2DB: data <= 32'b00000000000000000001000101100001;
				12'h2DC: data <= 32'b00000000000000000001000101110011;
				12'h2DD: data <= 32'b00000000000000000001000110000100;
				12'h2DE: data <= 32'b00000000000000000001000110010110;
				12'h2DF: data <= 32'b00000000000000000001000110101000;
				12'h2E0: data <= 32'b00000000000000000001000110111001;
				12'h2E1: data <= 32'b00000000000000000001000111001011;
				12'h2E2: data <= 32'b00000000000000000001000111011101;
				12'h2E3: data <= 32'b00000000000000000001000111101111;
				12'h2E4: data <= 32'b00000000000000000001001000000001;
				12'h2E5: data <= 32'b00000000000000000001001000010011;
				12'h2E6: data <= 32'b00000000000000000001001000100101;
				12'h2E7: data <= 32'b00000000000000000001001000110111;
				12'h2E8: data <= 32'b00000000000000000001001001001001;
				12'h2E9: data <= 32'b00000000000000000001001001011100;
				12'h2EA: data <= 32'b00000000000000000001001001101110;
				12'h2EB: data <= 32'b00000000000000000001001010000000;
				12'h2EC: data <= 32'b00000000000000000001001010010011;
				12'h2ED: data <= 32'b00000000000000000001001010100110;
				12'h2EE: data <= 32'b00000000000000000001001010111000;
				12'h2EF: data <= 32'b00000000000000000001001011001011;
				12'h2F0: data <= 32'b00000000000000000001001011011110;
				12'h2F1: data <= 32'b00000000000000000001001011110001;
				12'h2F2: data <= 32'b00000000000000000001001100000100;
				12'h2F3: data <= 32'b00000000000000000001001100010111;
				12'h2F4: data <= 32'b00000000000000000001001100101010;
				12'h2F5: data <= 32'b00000000000000000001001100111101;
				12'h2F6: data <= 32'b00000000000000000001001101010000;
				12'h2F7: data <= 32'b00000000000000000001001101100100;
				12'h2F8: data <= 32'b00000000000000000001001101110111;
				12'h2F9: data <= 32'b00000000000000000001001110001011;
				12'h2FA: data <= 32'b00000000000000000001001110011110;
				12'h2FB: data <= 32'b00000000000000000001001110110010;
				12'h2FC: data <= 32'b00000000000000000001001111000110;
				12'h2FD: data <= 32'b00000000000000000001001111011001;
				12'h2FE: data <= 32'b00000000000000000001001111101101;
				12'h2FF: data <= 32'b00000000000000000001010000000001;
				12'h300: data <= 32'b00000000000000000001010000010101;
				12'h301: data <= 32'b00000000000000000001010000101010;
				12'h302: data <= 32'b00000000000000000001010000111110;
				12'h303: data <= 32'b00000000000000000001010001010010;
				12'h304: data <= 32'b00000000000000000001010001100110;
				12'h305: data <= 32'b00000000000000000001010001111011;
				12'h306: data <= 32'b00000000000000000001010010001111;
				12'h307: data <= 32'b00000000000000000001010010100100;
				12'h308: data <= 32'b00000000000000000001010010111001;
				12'h309: data <= 32'b00000000000000000001010011001101;
				12'h30A: data <= 32'b00000000000000000001010011100010;
				12'h30B: data <= 32'b00000000000000000001010011110111;
				12'h30C: data <= 32'b00000000000000000001010100001100;
				12'h30D: data <= 32'b00000000000000000001010100100001;
				12'h30E: data <= 32'b00000000000000000001010100110110;
				12'h30F: data <= 32'b00000000000000000001010101001100;
				12'h310: data <= 32'b00000000000000000001010101100001;
				12'h311: data <= 32'b00000000000000000001010101110110;
				12'h312: data <= 32'b00000000000000000001010110001100;
				12'h313: data <= 32'b00000000000000000001010110100010;
				12'h314: data <= 32'b00000000000000000001010110110111;
				12'h315: data <= 32'b00000000000000000001010111001101;
				12'h316: data <= 32'b00000000000000000001010111100011;
				12'h317: data <= 32'b00000000000000000001010111111001;
				12'h318: data <= 32'b00000000000000000001011000001111;
				12'h319: data <= 32'b00000000000000000001011000100101;
				12'h31A: data <= 32'b00000000000000000001011000111011;
				12'h31B: data <= 32'b00000000000000000001011001010001;
				12'h31C: data <= 32'b00000000000000000001011001101000;
				12'h31D: data <= 32'b00000000000000000001011001111110;
				12'h31E: data <= 32'b00000000000000000001011010010101;
				12'h31F: data <= 32'b00000000000000000001011010101011;
				12'h320: data <= 32'b00000000000000000001011011000010;
				12'h321: data <= 32'b00000000000000000001011011011001;
				12'h322: data <= 32'b00000000000000000001011011110000;
				12'h323: data <= 32'b00000000000000000001011100000111;
				12'h324: data <= 32'b00000000000000000001011100011110;
				12'h325: data <= 32'b00000000000000000001011100110101;
				12'h326: data <= 32'b00000000000000000001011101001100;
				12'h327: data <= 32'b00000000000000000001011101100100;
				12'h328: data <= 32'b00000000000000000001011101111011;
				12'h329: data <= 32'b00000000000000000001011110010011;
				12'h32A: data <= 32'b00000000000000000001011110101010;
				12'h32B: data <= 32'b00000000000000000001011111000010;
				12'h32C: data <= 32'b00000000000000000001011111011010;
				12'h32D: data <= 32'b00000000000000000001011111110010;
				12'h32E: data <= 32'b00000000000000000001100000001010;
				12'h32F: data <= 32'b00000000000000000001100000100010;
				12'h330: data <= 32'b00000000000000000001100000111010;
				12'h331: data <= 32'b00000000000000000001100001010010;
				12'h332: data <= 32'b00000000000000000001100001101010;
				12'h333: data <= 32'b00000000000000000001100010000011;
				12'h334: data <= 32'b00000000000000000001100010011011;
				12'h335: data <= 32'b00000000000000000001100010110100;
				12'h336: data <= 32'b00000000000000000001100011001101;
				12'h337: data <= 32'b00000000000000000001100011100110;
				12'h338: data <= 32'b00000000000000000001100011111111;
				12'h339: data <= 32'b00000000000000000001100100011000;
				12'h33A: data <= 32'b00000000000000000001100100110001;
				12'h33B: data <= 32'b00000000000000000001100101001010;
				12'h33C: data <= 32'b00000000000000000001100101100011;
				12'h33D: data <= 32'b00000000000000000001100101111101;
				12'h33E: data <= 32'b00000000000000000001100110010110;
				12'h33F: data <= 32'b00000000000000000001100110110000;
				12'h340: data <= 32'b00000000000000000001100111001010;
				12'h341: data <= 32'b00000000000000000001100111100100;
				12'h342: data <= 32'b00000000000000000001100111111110;
				12'h343: data <= 32'b00000000000000000001101000011000;
				12'h344: data <= 32'b00000000000000000001101000110010;
				12'h345: data <= 32'b00000000000000000001101001001100;
				12'h346: data <= 32'b00000000000000000001101001100110;
				12'h347: data <= 32'b00000000000000000001101010000001;
				12'h348: data <= 32'b00000000000000000001101010011011;
				12'h349: data <= 32'b00000000000000000001101010110110;
				12'h34A: data <= 32'b00000000000000000001101011010001;
				12'h34B: data <= 32'b00000000000000000001101011101100;
				12'h34C: data <= 32'b00000000000000000001101100000111;
				12'h34D: data <= 32'b00000000000000000001101100100010;
				12'h34E: data <= 32'b00000000000000000001101100111101;
				12'h34F: data <= 32'b00000000000000000001101101011000;
				12'h350: data <= 32'b00000000000000000001101101110100;
				12'h351: data <= 32'b00000000000000000001101110001111;
				12'h352: data <= 32'b00000000000000000001101110101011;
				12'h353: data <= 32'b00000000000000000001101111000110;
				12'h354: data <= 32'b00000000000000000001101111100010;
				12'h355: data <= 32'b00000000000000000001101111111110;
				12'h356: data <= 32'b00000000000000000001110000011010;
				12'h357: data <= 32'b00000000000000000001110000110110;
				12'h358: data <= 32'b00000000000000000001110001010011;
				12'h359: data <= 32'b00000000000000000001110001101111;
				12'h35A: data <= 32'b00000000000000000001110010001100;
				12'h35B: data <= 32'b00000000000000000001110010101000;
				12'h35C: data <= 32'b00000000000000000001110011000101;
				12'h35D: data <= 32'b00000000000000000001110011100010;
				12'h35E: data <= 32'b00000000000000000001110011111111;
				12'h35F: data <= 32'b00000000000000000001110100011100;
				12'h360: data <= 32'b00000000000000000001110100111001;
				12'h361: data <= 32'b00000000000000000001110101010110;
				12'h362: data <= 32'b00000000000000000001110101110100;
				12'h363: data <= 32'b00000000000000000001110110010001;
				12'h364: data <= 32'b00000000000000000001110110101111;
				12'h365: data <= 32'b00000000000000000001110111001100;
				12'h366: data <= 32'b00000000000000000001110111101010;
				12'h367: data <= 32'b00000000000000000001111000001000;
				12'h368: data <= 32'b00000000000000000001111000100110;
				12'h369: data <= 32'b00000000000000000001111001000101;
				12'h36A: data <= 32'b00000000000000000001111001100011;
				12'h36B: data <= 32'b00000000000000000001111010000001;
				12'h36C: data <= 32'b00000000000000000001111010100000;
				12'h36D: data <= 32'b00000000000000000001111010111111;
				12'h36E: data <= 32'b00000000000000000001111011011101;
				12'h36F: data <= 32'b00000000000000000001111011111100;
				12'h370: data <= 32'b00000000000000000001111100011011;
				12'h371: data <= 32'b00000000000000000001111100111011;
				12'h372: data <= 32'b00000000000000000001111101011010;
				12'h373: data <= 32'b00000000000000000001111101111001;
				12'h374: data <= 32'b00000000000000000001111110011001;
				12'h375: data <= 32'b00000000000000000001111110111001;
				12'h376: data <= 32'b00000000000000000001111111011000;
				12'h377: data <= 32'b00000000000000000001111111111000;
				12'h378: data <= 32'b00000000000000000010000000011000;
				12'h379: data <= 32'b00000000000000000010000000111000;
				12'h37A: data <= 32'b00000000000000000010000001011001;
				12'h37B: data <= 32'b00000000000000000010000001111001;
				12'h37C: data <= 32'b00000000000000000010000010011010;
				12'h37D: data <= 32'b00000000000000000010000010111010;
				12'h37E: data <= 32'b00000000000000000010000011011011;
				12'h37F: data <= 32'b00000000000000000010000011111100;
				12'h380: data <= 32'b00000000000000000010000100011101;
				12'h381: data <= 32'b00000000000000000010000100111110;
				12'h382: data <= 32'b00000000000000000010000101100000;
				12'h383: data <= 32'b00000000000000000010000110000001;
				12'h384: data <= 32'b00000000000000000010000110100011;
				12'h385: data <= 32'b00000000000000000010000111000100;
				12'h386: data <= 32'b00000000000000000010000111100110;
				12'h387: data <= 32'b00000000000000000010001000001000;
				12'h388: data <= 32'b00000000000000000010001000101010;
				12'h389: data <= 32'b00000000000000000010001001001100;
				12'h38A: data <= 32'b00000000000000000010001001101111;
				12'h38B: data <= 32'b00000000000000000010001010010001;
				12'h38C: data <= 32'b00000000000000000010001010110100;
				12'h38D: data <= 32'b00000000000000000010001011010111;
				12'h38E: data <= 32'b00000000000000000010001011111010;
				12'h38F: data <= 32'b00000000000000000010001100011101;
				12'h390: data <= 32'b00000000000000000010001101000000;
				12'h391: data <= 32'b00000000000000000010001101100011;
				12'h392: data <= 32'b00000000000000000010001110000111;
				12'h393: data <= 32'b00000000000000000010001110101010;
				12'h394: data <= 32'b00000000000000000010001111001110;
				12'h395: data <= 32'b00000000000000000010001111110010;
				12'h396: data <= 32'b00000000000000000010010000010110;
				12'h397: data <= 32'b00000000000000000010010000111010;
				12'h398: data <= 32'b00000000000000000010010001011110;
				12'h399: data <= 32'b00000000000000000010010010000011;
				12'h39A: data <= 32'b00000000000000000010010010100111;
				12'h39B: data <= 32'b00000000000000000010010011001100;
				12'h39C: data <= 32'b00000000000000000010010011110001;
				12'h39D: data <= 32'b00000000000000000010010100010110;
				12'h39E: data <= 32'b00000000000000000010010100111011;
				12'h39F: data <= 32'b00000000000000000010010101100000;
				12'h3A0: data <= 32'b00000000000000000010010110000110;
				12'h3A1: data <= 32'b00000000000000000010010110101011;
				12'h3A2: data <= 32'b00000000000000000010010111010001;
				12'h3A3: data <= 32'b00000000000000000010010111110111;
				12'h3A4: data <= 32'b00000000000000000010011000011101;
				12'h3A5: data <= 32'b00000000000000000010011001000011;
				12'h3A6: data <= 32'b00000000000000000010011001101010;
				12'h3A7: data <= 32'b00000000000000000010011010010000;
				12'h3A8: data <= 32'b00000000000000000010011010110111;
				12'h3A9: data <= 32'b00000000000000000010011011011110;
				12'h3AA: data <= 32'b00000000000000000010011100000101;
				12'h3AB: data <= 32'b00000000000000000010011100101100;
				12'h3AC: data <= 32'b00000000000000000010011101010011;
				12'h3AD: data <= 32'b00000000000000000010011101111010;
				12'h3AE: data <= 32'b00000000000000000010011110100010;
				12'h3AF: data <= 32'b00000000000000000010011111001010;
				12'h3B0: data <= 32'b00000000000000000010011111110001;
				12'h3B1: data <= 32'b00000000000000000010100000011001;
				12'h3B2: data <= 32'b00000000000000000010100001000010;
				12'h3B3: data <= 32'b00000000000000000010100001101010;
				12'h3B4: data <= 32'b00000000000000000010100010010010;
				12'h3B5: data <= 32'b00000000000000000010100010111011;
				12'h3B6: data <= 32'b00000000000000000010100011100100;
				12'h3B7: data <= 32'b00000000000000000010100100001101;
				12'h3B8: data <= 32'b00000000000000000010100100110110;
				12'h3B9: data <= 32'b00000000000000000010100101011111;
				12'h3BA: data <= 32'b00000000000000000010100110001001;
				12'h3BB: data <= 32'b00000000000000000010100110110010;
				12'h3BC: data <= 32'b00000000000000000010100111011100;
				12'h3BD: data <= 32'b00000000000000000010101000000110;
				12'h3BE: data <= 32'b00000000000000000010101000110000;
				12'h3BF: data <= 32'b00000000000000000010101001011010;
				12'h3C0: data <= 32'b00000000000000000010101010000101;
				12'h3C1: data <= 32'b00000000000000000010101010110000;
				12'h3C2: data <= 32'b00000000000000000010101011011010;
				12'h3C3: data <= 32'b00000000000000000010101100000101;
				12'h3C4: data <= 32'b00000000000000000010101100110000;
				12'h3C5: data <= 32'b00000000000000000010101101011100;
				12'h3C6: data <= 32'b00000000000000000010101110000111;
				12'h3C7: data <= 32'b00000000000000000010101110110011;
				12'h3C8: data <= 32'b00000000000000000010101111011110;
				12'h3C9: data <= 32'b00000000000000000010110000001010;
				12'h3CA: data <= 32'b00000000000000000010110000110111;
				12'h3CB: data <= 32'b00000000000000000010110001100011;
				12'h3CC: data <= 32'b00000000000000000010110010001111;
				12'h3CD: data <= 32'b00000000000000000010110010111100;
				12'h3CE: data <= 32'b00000000000000000010110011101001;
				12'h3CF: data <= 32'b00000000000000000010110100010110;
				12'h3D0: data <= 32'b00000000000000000010110101000011;
				12'h3D1: data <= 32'b00000000000000000010110101110000;
				12'h3D2: data <= 32'b00000000000000000010110110011110;
				12'h3D3: data <= 32'b00000000000000000010110111001100;
				12'h3D4: data <= 32'b00000000000000000010110111111001;
				12'h3D5: data <= 32'b00000000000000000010111000100111;
				12'h3D6: data <= 32'b00000000000000000010111001010110;
				12'h3D7: data <= 32'b00000000000000000010111010000100;
				12'h3D8: data <= 32'b00000000000000000010111010110011;
				12'h3D9: data <= 32'b00000000000000000010111011100010;
				12'h3DA: data <= 32'b00000000000000000010111100010001;
				12'h3DB: data <= 32'b00000000000000000010111101000000;
				12'h3DC: data <= 32'b00000000000000000010111101101111;
				12'h3DD: data <= 32'b00000000000000000010111110011111;
				12'h3DE: data <= 32'b00000000000000000010111111001110;
				12'h3DF: data <= 32'b00000000000000000010111111111110;
				12'h3E0: data <= 32'b00000000000000000011000000101110;
				12'h3E1: data <= 32'b00000000000000000011000001011111;
				12'h3E2: data <= 32'b00000000000000000011000010001111;
				12'h3E3: data <= 32'b00000000000000000011000011000000;
				12'h3E4: data <= 32'b00000000000000000011000011110001;
				12'h3E5: data <= 32'b00000000000000000011000100100010;
				12'h3E6: data <= 32'b00000000000000000011000101010011;
				12'h3E7: data <= 32'b00000000000000000011000110000100;
				12'h3E8: data <= 32'b00000000000000000011000110110110;
				12'h3E9: data <= 32'b00000000000000000011000111101000;
				12'h3EA: data <= 32'b00000000000000000011001000011010;
				12'h3EB: data <= 32'b00000000000000000011001001001100;
				12'h3EC: data <= 32'b00000000000000000011001001111110;
				12'h3ED: data <= 32'b00000000000000000011001010110001;
				12'h3EE: data <= 32'b00000000000000000011001011100100;
				12'h3EF: data <= 32'b00000000000000000011001100010111;
				12'h3F0: data <= 32'b00000000000000000011001101001010;
				12'h3F1: data <= 32'b00000000000000000011001101111101;
				12'h3F2: data <= 32'b00000000000000000011001110110001;
				12'h3F3: data <= 32'b00000000000000000011001111100101;
				12'h3F4: data <= 32'b00000000000000000011010000011001;
				12'h3F5: data <= 32'b00000000000000000011010001001101;
				12'h3F6: data <= 32'b00000000000000000011010010000001;
				12'h3F7: data <= 32'b00000000000000000011010010110110;
				12'h3F8: data <= 32'b00000000000000000011010011101011;
				12'h3F9: data <= 32'b00000000000000000011010100100000;
				12'h3FA: data <= 32'b00000000000000000011010101010101;
				12'h3FB: data <= 32'b00000000000000000011010110001010;
				12'h3FC: data <= 32'b00000000000000000011010111000000;
				12'h3FD: data <= 32'b00000000000000000011010111110110;
				12'h3FE: data <= 32'b00000000000000000011011000101100;
				12'h3FF: data <= 32'b00000000000000000011011001100010;
				12'h400: data <= 32'b00000000000000000011011010011001;
				12'h401: data <= 32'b00000000000000000011011011001111;
				12'h402: data <= 32'b00000000000000000011011100000110;
				12'h403: data <= 32'b00000000000000000011011100111101;
				12'h404: data <= 32'b00000000000000000011011101110101;
				12'h405: data <= 32'b00000000000000000011011110101100;
				12'h406: data <= 32'b00000000000000000011011111100100;
				12'h407: data <= 32'b00000000000000000011100000011100;
				12'h408: data <= 32'b00000000000000000011100001010100;
				12'h409: data <= 32'b00000000000000000011100010001101;
				12'h40A: data <= 32'b00000000000000000011100011000101;
				12'h40B: data <= 32'b00000000000000000011100011111110;
				12'h40C: data <= 32'b00000000000000000011100100110111;
				12'h40D: data <= 32'b00000000000000000011100101110001;
				12'h40E: data <= 32'b00000000000000000011100110101010;
				12'h40F: data <= 32'b00000000000000000011100111100100;
				12'h410: data <= 32'b00000000000000000011101000011110;
				12'h411: data <= 32'b00000000000000000011101001011000;
				12'h412: data <= 32'b00000000000000000011101010010011;
				12'h413: data <= 32'b00000000000000000011101011001101;
				12'h414: data <= 32'b00000000000000000011101100001000;
				12'h415: data <= 32'b00000000000000000011101101000100;
				12'h416: data <= 32'b00000000000000000011101101111111;
				12'h417: data <= 32'b00000000000000000011101110111011;
				12'h418: data <= 32'b00000000000000000011101111110110;
				12'h419: data <= 32'b00000000000000000011110000110010;
				12'h41A: data <= 32'b00000000000000000011110001101111;
				12'h41B: data <= 32'b00000000000000000011110010101011;
				12'h41C: data <= 32'b00000000000000000011110011101000;
				12'h41D: data <= 32'b00000000000000000011110100100101;
				12'h41E: data <= 32'b00000000000000000011110101100010;
				12'h41F: data <= 32'b00000000000000000011110110100000;
				12'h420: data <= 32'b00000000000000000011110111011110;
				12'h421: data <= 32'b00000000000000000011111000011100;
				12'h422: data <= 32'b00000000000000000011111001011010;
				12'h423: data <= 32'b00000000000000000011111010011000;
				12'h424: data <= 32'b00000000000000000011111011010111;
				12'h425: data <= 32'b00000000000000000011111100010110;
				12'h426: data <= 32'b00000000000000000011111101010101;
				12'h427: data <= 32'b00000000000000000011111110010101;
				12'h428: data <= 32'b00000000000000000011111111010100;
				12'h429: data <= 32'b00000000000000000100000000010100;
				12'h42A: data <= 32'b00000000000000000100000001010101;
				12'h42B: data <= 32'b00000000000000000100000010010101;
				12'h42C: data <= 32'b00000000000000000100000011010110;
				12'h42D: data <= 32'b00000000000000000100000100010111;
				12'h42E: data <= 32'b00000000000000000100000101011000;
				12'h42F: data <= 32'b00000000000000000100000110011001;
				12'h430: data <= 32'b00000000000000000100000111011011;
				12'h431: data <= 32'b00000000000000000100001000011101;
				12'h432: data <= 32'b00000000000000000100001001011111;
				12'h433: data <= 32'b00000000000000000100001010100010;
				12'h434: data <= 32'b00000000000000000100001011100101;
				12'h435: data <= 32'b00000000000000000100001100101000;
				12'h436: data <= 32'b00000000000000000100001101101011;
				12'h437: data <= 32'b00000000000000000100001110101110;
				12'h438: data <= 32'b00000000000000000100001111110010;
				12'h439: data <= 32'b00000000000000000100010000110110;
				12'h43A: data <= 32'b00000000000000000100010001111011;
				12'h43B: data <= 32'b00000000000000000100010010111111;
				12'h43C: data <= 32'b00000000000000000100010100000100;
				12'h43D: data <= 32'b00000000000000000100010101001001;
				12'h43E: data <= 32'b00000000000000000100010110001111;
				12'h43F: data <= 32'b00000000000000000100010111010101;
				12'h440: data <= 32'b00000000000000000100011000011010;
				12'h441: data <= 32'b00000000000000000100011001100001;
				12'h442: data <= 32'b00000000000000000100011010100111;
				12'h443: data <= 32'b00000000000000000100011011101110;
				12'h444: data <= 32'b00000000000000000100011100110101;
				12'h445: data <= 32'b00000000000000000100011101111100;
				12'h446: data <= 32'b00000000000000000100011111000100;
				12'h447: data <= 32'b00000000000000000100100000001100;
				12'h448: data <= 32'b00000000000000000100100001010100;
				12'h449: data <= 32'b00000000000000000100100010011101;
				12'h44A: data <= 32'b00000000000000000100100011100101;
				12'h44B: data <= 32'b00000000000000000100100100101110;
				12'h44C: data <= 32'b00000000000000000100100101111000;
				12'h44D: data <= 32'b00000000000000000100100111000001;
				12'h44E: data <= 32'b00000000000000000100101000001011;
				12'h44F: data <= 32'b00000000000000000100101001010101;
				12'h450: data <= 32'b00000000000000000100101010100000;
				12'h451: data <= 32'b00000000000000000100101011101011;
				12'h452: data <= 32'b00000000000000000100101100110110;
				12'h453: data <= 32'b00000000000000000100101110000001;
				12'h454: data <= 32'b00000000000000000100101111001101;
				12'h455: data <= 32'b00000000000000000100110000011001;
				12'h456: data <= 32'b00000000000000000100110001100101;
				12'h457: data <= 32'b00000000000000000100110010110010;
				12'h458: data <= 32'b00000000000000000100110011111110;
				12'h459: data <= 32'b00000000000000000100110101001100;
				12'h45A: data <= 32'b00000000000000000100110110011001;
				12'h45B: data <= 32'b00000000000000000100110111100111;
				12'h45C: data <= 32'b00000000000000000100111000110101;
				12'h45D: data <= 32'b00000000000000000100111010000011;
				12'h45E: data <= 32'b00000000000000000100111011010010;
				12'h45F: data <= 32'b00000000000000000100111100100001;
				12'h460: data <= 32'b00000000000000000100111101110000;
				12'h461: data <= 32'b00000000000000000100111111000000;
				12'h462: data <= 32'b00000000000000000101000000010000;
				12'h463: data <= 32'b00000000000000000101000001100000;
				12'h464: data <= 32'b00000000000000000101000010110000;
				12'h465: data <= 32'b00000000000000000101000100000001;
				12'h466: data <= 32'b00000000000000000101000101010010;
				12'h467: data <= 32'b00000000000000000101000110100100;
				12'h468: data <= 32'b00000000000000000101000111110110;
				12'h469: data <= 32'b00000000000000000101001001001000;
				12'h46A: data <= 32'b00000000000000000101001010011010;
				12'h46B: data <= 32'b00000000000000000101001011101101;
				12'h46C: data <= 32'b00000000000000000101001101000000;
				12'h46D: data <= 32'b00000000000000000101001110010011;
				12'h46E: data <= 32'b00000000000000000101001111100111;
				12'h46F: data <= 32'b00000000000000000101010000111011;
				12'h470: data <= 32'b00000000000000000101010010010000;
				12'h471: data <= 32'b00000000000000000101010011100100;
				12'h472: data <= 32'b00000000000000000101010100111001;
				12'h473: data <= 32'b00000000000000000101010110001111;
				12'h474: data <= 32'b00000000000000000101010111100101;
				12'h475: data <= 32'b00000000000000000101011000111011;
				12'h476: data <= 32'b00000000000000000101011010010001;
				12'h477: data <= 32'b00000000000000000101011011101000;
				12'h478: data <= 32'b00000000000000000101011100111111;
				12'h479: data <= 32'b00000000000000000101011110010110;
				12'h47A: data <= 32'b00000000000000000101011111101110;
				12'h47B: data <= 32'b00000000000000000101100001000110;
				12'h47C: data <= 32'b00000000000000000101100010011111;
				12'h47D: data <= 32'b00000000000000000101100011110111;
				12'h47E: data <= 32'b00000000000000000101100101010001;
				12'h47F: data <= 32'b00000000000000000101100110101010;
				12'h480: data <= 32'b00000000000000000101101000000100;
				12'h481: data <= 32'b00000000000000000101101001011110;
				12'h482: data <= 32'b00000000000000000101101010111001;
				12'h483: data <= 32'b00000000000000000101101100010100;
				12'h484: data <= 32'b00000000000000000101101101101111;
				12'h485: data <= 32'b00000000000000000101101111001010;
				12'h486: data <= 32'b00000000000000000101110000100110;
				12'h487: data <= 32'b00000000000000000101110010000011;
				12'h488: data <= 32'b00000000000000000101110011011111;
				12'h489: data <= 32'b00000000000000000101110100111100;
				12'h48A: data <= 32'b00000000000000000101110110011010;
				12'h48B: data <= 32'b00000000000000000101110111111000;
				12'h48C: data <= 32'b00000000000000000101111001010110;
				12'h48D: data <= 32'b00000000000000000101111010110100;
				12'h48E: data <= 32'b00000000000000000101111100010011;
				12'h48F: data <= 32'b00000000000000000101111101110010;
				12'h490: data <= 32'b00000000000000000101111111010010;
				12'h491: data <= 32'b00000000000000000110000000110010;
				12'h492: data <= 32'b00000000000000000110000010010011;
				12'h493: data <= 32'b00000000000000000110000011110011;
				12'h494: data <= 32'b00000000000000000110000101010100;
				12'h495: data <= 32'b00000000000000000110000110110110;
				12'h496: data <= 32'b00000000000000000110001000011000;
				12'h497: data <= 32'b00000000000000000110001001111010;
				12'h498: data <= 32'b00000000000000000110001011011101;
				12'h499: data <= 32'b00000000000000000110001101000000;
				12'h49A: data <= 32'b00000000000000000110001110100011;
				12'h49B: data <= 32'b00000000000000000110010000000111;
				12'h49C: data <= 32'b00000000000000000110010001101011;
				12'h49D: data <= 32'b00000000000000000110010011010000;
				12'h49E: data <= 32'b00000000000000000110010100110101;
				12'h49F: data <= 32'b00000000000000000110010110011010;
				12'h4A0: data <= 32'b00000000000000000110011000000000;
				12'h4A1: data <= 32'b00000000000000000110011001100110;
				12'h4A2: data <= 32'b00000000000000000110011011001101;
				12'h4A3: data <= 32'b00000000000000000110011100110100;
				12'h4A4: data <= 32'b00000000000000000110011110011011;
				12'h4A5: data <= 32'b00000000000000000110100000000011;
				12'h4A6: data <= 32'b00000000000000000110100001101011;
				12'h4A7: data <= 32'b00000000000000000110100011010100;
				12'h4A8: data <= 32'b00000000000000000110100100111101;
				12'h4A9: data <= 32'b00000000000000000110100110100111;
				12'h4AA: data <= 32'b00000000000000000110101000010000;
				12'h4AB: data <= 32'b00000000000000000110101001111011;
				12'h4AC: data <= 32'b00000000000000000110101011100101;
				12'h4AD: data <= 32'b00000000000000000110101101010000;
				12'h4AE: data <= 32'b00000000000000000110101110111100;
				12'h4AF: data <= 32'b00000000000000000110110000101000;
				12'h4B0: data <= 32'b00000000000000000110110010010100;
				12'h4B1: data <= 32'b00000000000000000110110100000001;
				12'h4B2: data <= 32'b00000000000000000110110101101110;
				12'h4B3: data <= 32'b00000000000000000110110111011100;
				12'h4B4: data <= 32'b00000000000000000110111001001010;
				12'h4B5: data <= 32'b00000000000000000110111010111001;
				12'h4B6: data <= 32'b00000000000000000110111100101000;
				12'h4B7: data <= 32'b00000000000000000110111110010111;
				12'h4B8: data <= 32'b00000000000000000111000000000111;
				12'h4B9: data <= 32'b00000000000000000111000001110111;
				12'h4BA: data <= 32'b00000000000000000111000011101000;
				12'h4BB: data <= 32'b00000000000000000111000101011001;
				12'h4BC: data <= 32'b00000000000000000111000111001010;
				12'h4BD: data <= 32'b00000000000000000111001000111100;
				12'h4BE: data <= 32'b00000000000000000111001010101111;
				12'h4BF: data <= 32'b00000000000000000111001100100010;
				12'h4C0: data <= 32'b00000000000000000111001110010101;
				12'h4C1: data <= 32'b00000000000000000111010000001001;
				12'h4C2: data <= 32'b00000000000000000111010001111101;
				12'h4C3: data <= 32'b00000000000000000111010011110010;
				12'h4C4: data <= 32'b00000000000000000111010101100111;
				12'h4C5: data <= 32'b00000000000000000111010111011101;
				12'h4C6: data <= 32'b00000000000000000111011001010011;
				12'h4C7: data <= 32'b00000000000000000111011011001001;
				12'h4C8: data <= 32'b00000000000000000111011101000000;
				12'h4C9: data <= 32'b00000000000000000111011110111000;
				12'h4CA: data <= 32'b00000000000000000111100000110000;
				12'h4CB: data <= 32'b00000000000000000111100010101000;
				12'h4CC: data <= 32'b00000000000000000111100100100001;
				12'h4CD: data <= 32'b00000000000000000111100110011010;
				12'h4CE: data <= 32'b00000000000000000111101000010100;
				12'h4CF: data <= 32'b00000000000000000111101010001111;
				12'h4D0: data <= 32'b00000000000000000111101100001001;
				12'h4D1: data <= 32'b00000000000000000111101110000101;
				12'h4D2: data <= 32'b00000000000000000111110000000000;
				12'h4D3: data <= 32'b00000000000000000111110001111101;
				12'h4D4: data <= 32'b00000000000000000111110011111001;
				12'h4D5: data <= 32'b00000000000000000111110101110111;
				12'h4D6: data <= 32'b00000000000000000111110111110100;
				12'h4D7: data <= 32'b00000000000000000111111001110011;
				12'h4D8: data <= 32'b00000000000000000111111011110001;
				12'h4D9: data <= 32'b00000000000000000111111101110000;
				12'h4DA: data <= 32'b00000000000000000111111111110000;
				12'h4DB: data <= 32'b00000000000000001000000001110000;
				12'h4DC: data <= 32'b00000000000000001000000011110001;
				12'h4DD: data <= 32'b00000000000000001000000101110010;
				12'h4DE: data <= 32'b00000000000000001000000111110100;
				12'h4DF: data <= 32'b00000000000000001000001001110110;
				12'h4E0: data <= 32'b00000000000000001000001011111001;
				12'h4E1: data <= 32'b00000000000000001000001101111100;
				12'h4E2: data <= 32'b00000000000000001000010000000000;
				12'h4E3: data <= 32'b00000000000000001000010010000100;
				12'h4E4: data <= 32'b00000000000000001000010100001001;
				12'h4E5: data <= 32'b00000000000000001000010110001110;
				12'h4E6: data <= 32'b00000000000000001000011000010100;
				12'h4E7: data <= 32'b00000000000000001000011010011010;
				12'h4E8: data <= 32'b00000000000000001000011100100001;
				12'h4E9: data <= 32'b00000000000000001000011110101001;
				12'h4EA: data <= 32'b00000000000000001000100000110001;
				12'h4EB: data <= 32'b00000000000000001000100010111001;
				12'h4EC: data <= 32'b00000000000000001000100101000010;
				12'h4ED: data <= 32'b00000000000000001000100111001100;
				12'h4EE: data <= 32'b00000000000000001000101001010110;
				12'h4EF: data <= 32'b00000000000000001000101011100000;
				12'h4F0: data <= 32'b00000000000000001000101101101011;
				12'h4F1: data <= 32'b00000000000000001000101111110111;
				12'h4F2: data <= 32'b00000000000000001000110010000011;
				12'h4F3: data <= 32'b00000000000000001000110100010000;
				12'h4F4: data <= 32'b00000000000000001000110110011101;
				12'h4F5: data <= 32'b00000000000000001000111000101011;
				12'h4F6: data <= 32'b00000000000000001000111010111010;
				12'h4F7: data <= 32'b00000000000000001000111101001001;
				12'h4F8: data <= 32'b00000000000000001000111111011000;
				12'h4F9: data <= 32'b00000000000000001001000001101000;
				12'h4FA: data <= 32'b00000000000000001001000011111001;
				12'h4FB: data <= 32'b00000000000000001001000110001010;
				12'h4FC: data <= 32'b00000000000000001001001000011100;
				12'h4FD: data <= 32'b00000000000000001001001010101111;
				12'h4FE: data <= 32'b00000000000000001001001101000010;
				12'h4FF: data <= 32'b00000000000000001001001111010101;
				12'h500: data <= 32'b00000000000000001001010001101001;
				12'h501: data <= 32'b00000000000000001001010011111110;
				12'h502: data <= 32'b00000000000000001001010110010011;
				12'h503: data <= 32'b00000000000000001001011000101001;
				12'h504: data <= 32'b00000000000000001001011011000000;
				12'h505: data <= 32'b00000000000000001001011101010111;
				12'h506: data <= 32'b00000000000000001001011111101110;
				12'h507: data <= 32'b00000000000000001001100010000110;
				12'h508: data <= 32'b00000000000000001001100100011111;
				12'h509: data <= 32'b00000000000000001001100110111001;
				12'h50A: data <= 32'b00000000000000001001101001010011;
				12'h50B: data <= 32'b00000000000000001001101011101101;
				12'h50C: data <= 32'b00000000000000001001101110001001;
				12'h50D: data <= 32'b00000000000000001001110000100100;
				12'h50E: data <= 32'b00000000000000001001110011000001;
				12'h50F: data <= 32'b00000000000000001001110101011110;
				12'h510: data <= 32'b00000000000000001001110111111100;
				12'h511: data <= 32'b00000000000000001001111010011010;
				12'h512: data <= 32'b00000000000000001001111100111001;
				12'h513: data <= 32'b00000000000000001001111111011000;
				12'h514: data <= 32'b00000000000000001010000001111001;
				12'h515: data <= 32'b00000000000000001010000100011001;
				12'h516: data <= 32'b00000000000000001010000110111011;
				12'h517: data <= 32'b00000000000000001010001001011101;
				12'h518: data <= 32'b00000000000000001010001011111111;
				12'h519: data <= 32'b00000000000000001010001110100011;
				12'h51A: data <= 32'b00000000000000001010010001000111;
				12'h51B: data <= 32'b00000000000000001010010011101011;
				12'h51C: data <= 32'b00000000000000001010010110010001;
				12'h51D: data <= 32'b00000000000000001010011000110111;
				12'h51E: data <= 32'b00000000000000001010011011011101;
				12'h51F: data <= 32'b00000000000000001010011110000100;
				12'h520: data <= 32'b00000000000000001010100000101100;
				12'h521: data <= 32'b00000000000000001010100011010101;
				12'h522: data <= 32'b00000000000000001010100101111110;
				12'h523: data <= 32'b00000000000000001010101000101000;
				12'h524: data <= 32'b00000000000000001010101011010010;
				12'h525: data <= 32'b00000000000000001010101101111101;
				12'h526: data <= 32'b00000000000000001010110000101001;
				12'h527: data <= 32'b00000000000000001010110011010110;
				12'h528: data <= 32'b00000000000000001010110110000011;
				12'h529: data <= 32'b00000000000000001010111000110001;
				12'h52A: data <= 32'b00000000000000001010111011011111;
				12'h52B: data <= 32'b00000000000000001010111110001110;
				12'h52C: data <= 32'b00000000000000001011000000111110;
				12'h52D: data <= 32'b00000000000000001011000011101111;
				12'h52E: data <= 32'b00000000000000001011000110100000;
				12'h52F: data <= 32'b00000000000000001011001001010010;
				12'h530: data <= 32'b00000000000000001011001100000101;
				12'h531: data <= 32'b00000000000000001011001110111000;
				12'h532: data <= 32'b00000000000000001011010001101100;
				12'h533: data <= 32'b00000000000000001011010100100001;
				12'h534: data <= 32'b00000000000000001011010111010110;
				12'h535: data <= 32'b00000000000000001011011010001101;
				12'h536: data <= 32'b00000000000000001011011101000100;
				12'h537: data <= 32'b00000000000000001011011111111011;
				12'h538: data <= 32'b00000000000000001011100010110100;
				12'h539: data <= 32'b00000000000000001011100101101101;
				12'h53A: data <= 32'b00000000000000001011101000100110;
				12'h53B: data <= 32'b00000000000000001011101011100001;
				12'h53C: data <= 32'b00000000000000001011101110011100;
				12'h53D: data <= 32'b00000000000000001011110001011000;
				12'h53E: data <= 32'b00000000000000001011110100010101;
				12'h53F: data <= 32'b00000000000000001011110111010010;
				12'h540: data <= 32'b00000000000000001011111010010000;
				12'h541: data <= 32'b00000000000000001011111101001111;
				12'h542: data <= 32'b00000000000000001100000000001111;
				12'h543: data <= 32'b00000000000000001100000011010000;
				12'h544: data <= 32'b00000000000000001100000110010001;
				12'h545: data <= 32'b00000000000000001100001001010011;
				12'h546: data <= 32'b00000000000000001100001100010101;
				12'h547: data <= 32'b00000000000000001100001111011001;
				12'h548: data <= 32'b00000000000000001100010010011101;
				12'h549: data <= 32'b00000000000000001100010101100010;
				12'h54A: data <= 32'b00000000000000001100011000101000;
				12'h54B: data <= 32'b00000000000000001100011011101110;
				12'h54C: data <= 32'b00000000000000001100011110110110;
				12'h54D: data <= 32'b00000000000000001100100001111110;
				12'h54E: data <= 32'b00000000000000001100100101000111;
				12'h54F: data <= 32'b00000000000000001100101000010000;
				12'h550: data <= 32'b00000000000000001100101011011011;
				12'h551: data <= 32'b00000000000000001100101110100110;
				12'h552: data <= 32'b00000000000000001100110001110010;
				12'h553: data <= 32'b00000000000000001100110100111111;
				12'h554: data <= 32'b00000000000000001100111000001101;
				12'h555: data <= 32'b00000000000000001100111011011011;
				12'h556: data <= 32'b00000000000000001100111110101010;
				12'h557: data <= 32'b00000000000000001101000001111010;
				12'h558: data <= 32'b00000000000000001101000101001011;
				12'h559: data <= 32'b00000000000000001101001000011101;
				12'h55A: data <= 32'b00000000000000001101001011110000;
				12'h55B: data <= 32'b00000000000000001101001111000011;
				12'h55C: data <= 32'b00000000000000001101010010010111;
				12'h55D: data <= 32'b00000000000000001101010101101100;
				12'h55E: data <= 32'b00000000000000001101011001000010;
				12'h55F: data <= 32'b00000000000000001101011100011001;
				12'h560: data <= 32'b00000000000000001101011111110000;
				12'h561: data <= 32'b00000000000000001101100011001000;
				12'h562: data <= 32'b00000000000000001101100110100010;
				12'h563: data <= 32'b00000000000000001101101001111100;
				12'h564: data <= 32'b00000000000000001101101101010111;
				12'h565: data <= 32'b00000000000000001101110000110010;
				12'h566: data <= 32'b00000000000000001101110100001111;
				12'h567: data <= 32'b00000000000000001101110111101101;
				12'h568: data <= 32'b00000000000000001101111011001011;
				12'h569: data <= 32'b00000000000000001101111110101010;
				12'h56A: data <= 32'b00000000000000001110000010001010;
				12'h56B: data <= 32'b00000000000000001110000101101011;
				12'h56C: data <= 32'b00000000000000001110001001001101;
				12'h56D: data <= 32'b00000000000000001110001100110000;
				12'h56E: data <= 32'b00000000000000001110010000010011;
				12'h56F: data <= 32'b00000000000000001110010011111000;
				12'h570: data <= 32'b00000000000000001110010111011101;
				12'h571: data <= 32'b00000000000000001110011011000100;
				12'h572: data <= 32'b00000000000000001110011110101011;
				12'h573: data <= 32'b00000000000000001110100010010011;
				12'h574: data <= 32'b00000000000000001110100101111100;
				12'h575: data <= 32'b00000000000000001110101001100110;
				12'h576: data <= 32'b00000000000000001110101101010001;
				12'h577: data <= 32'b00000000000000001110110000111101;
				12'h578: data <= 32'b00000000000000001110110100101001;
				12'h579: data <= 32'b00000000000000001110111000010111;
				12'h57A: data <= 32'b00000000000000001110111100000110;
				12'h57B: data <= 32'b00000000000000001110111111110101;
				12'h57C: data <= 32'b00000000000000001111000011100101;
				12'h57D: data <= 32'b00000000000000001111000111010111;
				12'h57E: data <= 32'b00000000000000001111001011001001;
				12'h57F: data <= 32'b00000000000000001111001110111100;
				12'h580: data <= 32'b00000000000000001111010010110001;
				12'h581: data <= 32'b00000000000000001111010110100110;
				12'h582: data <= 32'b00000000000000001111011010011100;
				12'h583: data <= 32'b00000000000000001111011110010011;
				12'h584: data <= 32'b00000000000000001111100010001011;
				12'h585: data <= 32'b00000000000000001111100110000100;
				12'h586: data <= 32'b00000000000000001111101001111110;
				12'h587: data <= 32'b00000000000000001111101101111001;
				12'h588: data <= 32'b00000000000000001111110001110101;
				12'h589: data <= 32'b00000000000000001111110101110010;
				12'h58A: data <= 32'b00000000000000001111111001110000;
				12'h58B: data <= 32'b00000000000000001111111101101111;
				12'h58C: data <= 32'b00000000000000010000000001101111;
				12'h58D: data <= 32'b00000000000000010000000101110000;
				12'h58E: data <= 32'b00000000000000010000001001110010;
				12'h58F: data <= 32'b00000000000000010000001101110101;
				12'h590: data <= 32'b00000000000000010000010001111001;
				12'h591: data <= 32'b00000000000000010000010101111110;
				12'h592: data <= 32'b00000000000000010000011010000100;
				12'h593: data <= 32'b00000000000000010000011110001011;
				12'h594: data <= 32'b00000000000000010000100010010011;
				12'h595: data <= 32'b00000000000000010000100110011100;
				12'h596: data <= 32'b00000000000000010000101010100110;
				12'h597: data <= 32'b00000000000000010000101110110001;
				12'h598: data <= 32'b00000000000000010000110010111101;
				12'h599: data <= 32'b00000000000000010000110111001011;
				12'h59A: data <= 32'b00000000000000010000111011011001;
				12'h59B: data <= 32'b00000000000000010000111111101000;
				12'h59C: data <= 32'b00000000000000010001000011111001;
				12'h59D: data <= 32'b00000000000000010001001000001010;
				12'h59E: data <= 32'b00000000000000010001001100011101;
				12'h59F: data <= 32'b00000000000000010001010000110000;
				12'h5A0: data <= 32'b00000000000000010001010101000101;
				12'h5A1: data <= 32'b00000000000000010001011001011011;
				12'h5A2: data <= 32'b00000000000000010001011101110010;
				12'h5A3: data <= 32'b00000000000000010001100010001010;
				12'h5A4: data <= 32'b00000000000000010001100110100011;
				12'h5A5: data <= 32'b00000000000000010001101010111101;
				12'h5A6: data <= 32'b00000000000000010001101111011000;
				12'h5A7: data <= 32'b00000000000000010001110011110101;
				12'h5A8: data <= 32'b00000000000000010001111000010010;
				12'h5A9: data <= 32'b00000000000000010001111100110001;
				12'h5AA: data <= 32'b00000000000000010010000001010001;
				12'h5AB: data <= 32'b00000000000000010010000101110010;
				12'h5AC: data <= 32'b00000000000000010010001010010100;
				12'h5AD: data <= 32'b00000000000000010010001110110111;
				12'h5AE: data <= 32'b00000000000000010010010011011011;
				12'h5AF: data <= 32'b00000000000000010010011000000001;
				12'h5B0: data <= 32'b00000000000000010010011100100111;
				12'h5B1: data <= 32'b00000000000000010010100001001111;
				12'h5B2: data <= 32'b00000000000000010010100101111000;
				12'h5B3: data <= 32'b00000000000000010010101010100010;
				12'h5B4: data <= 32'b00000000000000010010101111001101;
				12'h5B5: data <= 32'b00000000000000010010110011111001;
				12'h5B6: data <= 32'b00000000000000010010111000100111;
				12'h5B7: data <= 32'b00000000000000010010111101010110;
				12'h5B8: data <= 32'b00000000000000010011000010000110;
				12'h5B9: data <= 32'b00000000000000010011000110110111;
				12'h5BA: data <= 32'b00000000000000010011001011101001;
				12'h5BB: data <= 32'b00000000000000010011010000011101;
				12'h5BC: data <= 32'b00000000000000010011010101010001;
				12'h5BD: data <= 32'b00000000000000010011011010000111;
				12'h5BE: data <= 32'b00000000000000010011011110111110;
				12'h5BF: data <= 32'b00000000000000010011100011110111;
				12'h5C0: data <= 32'b00000000000000010011101000110000;
				12'h5C1: data <= 32'b00000000000000010011101101101011;
				12'h5C2: data <= 32'b00000000000000010011110010100111;
				12'h5C3: data <= 32'b00000000000000010011110111100100;
				12'h5C4: data <= 32'b00000000000000010011111100100011;
				12'h5C5: data <= 32'b00000000000000010100000001100011;
				12'h5C6: data <= 32'b00000000000000010100000110100100;
				12'h5C7: data <= 32'b00000000000000010100001011100110;
				12'h5C8: data <= 32'b00000000000000010100010000101010;
				12'h5C9: data <= 32'b00000000000000010100010101101110;
				12'h5CA: data <= 32'b00000000000000010100011010110100;
				12'h5CB: data <= 32'b00000000000000010100011111111100;
				12'h5CC: data <= 32'b00000000000000010100100101000100;
				12'h5CD: data <= 32'b00000000000000010100101010001110;
				12'h5CE: data <= 32'b00000000000000010100101111011001;
				12'h5CF: data <= 32'b00000000000000010100110100100110;
				12'h5D0: data <= 32'b00000000000000010100111001110100;
				12'h5D1: data <= 32'b00000000000000010100111111000011;
				12'h5D2: data <= 32'b00000000000000010101000100010011;
				12'h5D3: data <= 32'b00000000000000010101001001100101;
				12'h5D4: data <= 32'b00000000000000010101001110111000;
				12'h5D5: data <= 32'b00000000000000010101010100001100;
				12'h5D6: data <= 32'b00000000000000010101011001100010;
				12'h5D7: data <= 32'b00000000000000010101011110111001;
				12'h5D8: data <= 32'b00000000000000010101100100010010;
				12'h5D9: data <= 32'b00000000000000010101101001101011;
				12'h5DA: data <= 32'b00000000000000010101101111000111;
				12'h5DB: data <= 32'b00000000000000010101110100100011;
				12'h5DC: data <= 32'b00000000000000010101111010000001;
				12'h5DD: data <= 32'b00000000000000010101111111100000;
				12'h5DE: data <= 32'b00000000000000010110000101000001;
				12'h5DF: data <= 32'b00000000000000010110001010100010;
				12'h5E0: data <= 32'b00000000000000010110010000000110;
				12'h5E1: data <= 32'b00000000000000010110010101101011;
				12'h5E2: data <= 32'b00000000000000010110011011010001;
				12'h5E3: data <= 32'b00000000000000010110100000111000;
				12'h5E4: data <= 32'b00000000000000010110100110100001;
				12'h5E5: data <= 32'b00000000000000010110101100001011;
				12'h5E6: data <= 32'b00000000000000010110110001110111;
				12'h5E7: data <= 32'b00000000000000010110110111100100;
				12'h5E8: data <= 32'b00000000000000010110111101010011;
				12'h5E9: data <= 32'b00000000000000010111000011000011;
				12'h5EA: data <= 32'b00000000000000010111001000110101;
				12'h5EB: data <= 32'b00000000000000010111001110100111;
				12'h5EC: data <= 32'b00000000000000010111010100011100;
				12'h5ED: data <= 32'b00000000000000010111011010010010;
				12'h5EE: data <= 32'b00000000000000010111100000001001;
				12'h5EF: data <= 32'b00000000000000010111100110000010;
				12'h5F0: data <= 32'b00000000000000010111101011111100;
				12'h5F1: data <= 32'b00000000000000010111110001111000;
				12'h5F2: data <= 32'b00000000000000010111110111110101;
				12'h5F3: data <= 32'b00000000000000010111111101110100;
				12'h5F4: data <= 32'b00000000000000011000000011110100;
				12'h5F5: data <= 32'b00000000000000011000001001110110;
				12'h5F6: data <= 32'b00000000000000011000001111111001;
				12'h5F7: data <= 32'b00000000000000011000010101111101;
				12'h5F8: data <= 32'b00000000000000011000011100000100;
				12'h5F9: data <= 32'b00000000000000011000100010001100;
				12'h5FA: data <= 32'b00000000000000011000101000010101;
				12'h5FB: data <= 32'b00000000000000011000101110100000;
				12'h5FC: data <= 32'b00000000000000011000110100101100;
				12'h5FD: data <= 32'b00000000000000011000111010111010;
				12'h5FE: data <= 32'b00000000000000011001000001001010;
				12'h5FF: data <= 32'b00000000000000011001000111011011;
				12'h600: data <= 32'b00000000000000011001001101101101;
				12'h601: data <= 32'b00000000000000011001010100000001;
				12'h602: data <= 32'b00000000000000011001011010010111;
				12'h603: data <= 32'b00000000000000011001100000101111;
				12'h604: data <= 32'b00000000000000011001100111001000;
				12'h605: data <= 32'b00000000000000011001101101100010;
				12'h606: data <= 32'b00000000000000011001110011111110;
				12'h607: data <= 32'b00000000000000011001111010011100;
				12'h608: data <= 32'b00000000000000011010000000111100;
				12'h609: data <= 32'b00000000000000011010000111011101;
				12'h60A: data <= 32'b00000000000000011010001101111111;
				12'h60B: data <= 32'b00000000000000011010010100100100;
				12'h60C: data <= 32'b00000000000000011010011011001010;
				12'h60D: data <= 32'b00000000000000011010100001110001;
				12'h60E: data <= 32'b00000000000000011010101000011011;
				12'h60F: data <= 32'b00000000000000011010101111000110;
				12'h610: data <= 32'b00000000000000011010110101110010;
				12'h611: data <= 32'b00000000000000011010111100100000;
				12'h612: data <= 32'b00000000000000011011000011010000;
				12'h613: data <= 32'b00000000000000011011001010000010;
				12'h614: data <= 32'b00000000000000011011010000110101;
				12'h615: data <= 32'b00000000000000011011010111101010;
				12'h616: data <= 32'b00000000000000011011011110100001;
				12'h617: data <= 32'b00000000000000011011100101011010;
				12'h618: data <= 32'b00000000000000011011101100010100;
				12'h619: data <= 32'b00000000000000011011110011010000;
				12'h61A: data <= 32'b00000000000000011011111010001110;
				12'h61B: data <= 32'b00000000000000011100000001001101;
				12'h61C: data <= 32'b00000000000000011100001000001110;
				12'h61D: data <= 32'b00000000000000011100001111010001;
				12'h61E: data <= 32'b00000000000000011100010110010110;
				12'h61F: data <= 32'b00000000000000011100011101011100;
				12'h620: data <= 32'b00000000000000011100100100100101;
				12'h621: data <= 32'b00000000000000011100101011101111;
				12'h622: data <= 32'b00000000000000011100110010111010;
				12'h623: data <= 32'b00000000000000011100111010001000;
				12'h624: data <= 32'b00000000000000011101000001010111;
				12'h625: data <= 32'b00000000000000011101001000101001;
				12'h626: data <= 32'b00000000000000011101001111111100;
				12'h627: data <= 32'b00000000000000011101010111010001;
				12'h628: data <= 32'b00000000000000011101011110100111;
				12'h629: data <= 32'b00000000000000011101100110000000;
				12'h62A: data <= 32'b00000000000000011101101101011010;
				12'h62B: data <= 32'b00000000000000011101110100110111;
				12'h62C: data <= 32'b00000000000000011101111100010101;
				12'h62D: data <= 32'b00000000000000011110000011110101;
				12'h62E: data <= 32'b00000000000000011110001011010111;
				12'h62F: data <= 32'b00000000000000011110010010111011;
				12'h630: data <= 32'b00000000000000011110011010100000;
				12'h631: data <= 32'b00000000000000011110100010001000;
				12'h632: data <= 32'b00000000000000011110101001110001;
				12'h633: data <= 32'b00000000000000011110110001011101;
				12'h634: data <= 32'b00000000000000011110111001001010;
				12'h635: data <= 32'b00000000000000011111000000111001;
				12'h636: data <= 32'b00000000000000011111001000101011;
				12'h637: data <= 32'b00000000000000011111010000011110;
				12'h638: data <= 32'b00000000000000011111011000010011;
				12'h639: data <= 32'b00000000000000011111100000001010;
				12'h63A: data <= 32'b00000000000000011111101000000011;
				12'h63B: data <= 32'b00000000000000011111101111111110;
				12'h63C: data <= 32'b00000000000000011111110111111011;
				12'h63D: data <= 32'b00000000000000011111111111111010;
				12'h63E: data <= 32'b00000000000000100000000111111011;
				12'h63F: data <= 32'b00000000000000100000001111111110;
				12'h640: data <= 32'b00000000000000100000011000000011;
				12'h641: data <= 32'b00000000000000100000100000001010;
				12'h642: data <= 32'b00000000000000100000101000010011;
				12'h643: data <= 32'b00000000000000100000110000011110;
				12'h644: data <= 32'b00000000000000100000111000101011;
				12'h645: data <= 32'b00000000000000100001000000111010;
				12'h646: data <= 32'b00000000000000100001001001001100;
				12'h647: data <= 32'b00000000000000100001010001011111;
				12'h648: data <= 32'b00000000000000100001011001110100;
				12'h649: data <= 32'b00000000000000100001100010001100;
				12'h64A: data <= 32'b00000000000000100001101010100101;
				12'h64B: data <= 32'b00000000000000100001110011000001;
				12'h64C: data <= 32'b00000000000000100001111011011111;
				12'h64D: data <= 32'b00000000000000100010000011111111;
				12'h64E: data <= 32'b00000000000000100010001100100001;
				12'h64F: data <= 32'b00000000000000100010010101000101;
				12'h650: data <= 32'b00000000000000100010011101101011;
				12'h651: data <= 32'b00000000000000100010100110010100;
				12'h652: data <= 32'b00000000000000100010101110111111;
				12'h653: data <= 32'b00000000000000100010110111101011;
				12'h654: data <= 32'b00000000000000100011000000011010;
				12'h655: data <= 32'b00000000000000100011001001001100;
				12'h656: data <= 32'b00000000000000100011010001111111;
				12'h657: data <= 32'b00000000000000100011011010110101;
				12'h658: data <= 32'b00000000000000100011100011101101;
				12'h659: data <= 32'b00000000000000100011101100100111;
				12'h65A: data <= 32'b00000000000000100011110101100011;
				12'h65B: data <= 32'b00000000000000100011111110100001;
				12'h65C: data <= 32'b00000000000000100100000111100010;
				12'h65D: data <= 32'b00000000000000100100010000100101;
				12'h65E: data <= 32'b00000000000000100100011001101010;
				12'h65F: data <= 32'b00000000000000100100100010110010;
				12'h660: data <= 32'b00000000000000100100101011111100;
				12'h661: data <= 32'b00000000000000100100110101001000;
				12'h662: data <= 32'b00000000000000100100111110010110;
				12'h663: data <= 32'b00000000000000100101000111100111;
				12'h664: data <= 32'b00000000000000100101010000111010;
				12'h665: data <= 32'b00000000000000100101011010010000;
				12'h666: data <= 32'b00000000000000100101100011100111;
				12'h667: data <= 32'b00000000000000100101101101000001;
				12'h668: data <= 32'b00000000000000100101110110011110;
				12'h669: data <= 32'b00000000000000100101111111111101;
				12'h66A: data <= 32'b00000000000000100110001001011110;
				12'h66B: data <= 32'b00000000000000100110010011000001;
				12'h66C: data <= 32'b00000000000000100110011100100111;
				12'h66D: data <= 32'b00000000000000100110100110010000;
				12'h66E: data <= 32'b00000000000000100110101111111010;
				12'h66F: data <= 32'b00000000000000100110111001101000;
				12'h670: data <= 32'b00000000000000100111000011010111;
				12'h671: data <= 32'b00000000000000100111001101001001;
				12'h672: data <= 32'b00000000000000100111010110111110;
				12'h673: data <= 32'b00000000000000100111100000110101;
				12'h674: data <= 32'b00000000000000100111101010101110;
				12'h675: data <= 32'b00000000000000100111110100101010;
				12'h676: data <= 32'b00000000000000100111111110101001;
				12'h677: data <= 32'b00000000000000101000001000101001;
				12'h678: data <= 32'b00000000000000101000010010101101;
				12'h679: data <= 32'b00000000000000101000011100110011;
				12'h67A: data <= 32'b00000000000000101000100110111011;
				12'h67B: data <= 32'b00000000000000101000110001000110;
				12'h67C: data <= 32'b00000000000000101000111011010100;
				12'h67D: data <= 32'b00000000000000101001000101100100;
				12'h67E: data <= 32'b00000000000000101001001111110111;
				12'h67F: data <= 32'b00000000000000101001011010001100;
				12'h680: data <= 32'b00000000000000101001100100100100;
				12'h681: data <= 32'b00000000000000101001101110111110;
				12'h682: data <= 32'b00000000000000101001111001011011;
				12'h683: data <= 32'b00000000000000101010000011111011;
				12'h684: data <= 32'b00000000000000101010001110011101;
				12'h685: data <= 32'b00000000000000101010011001000010;
				12'h686: data <= 32'b00000000000000101010100011101010;
				12'h687: data <= 32'b00000000000000101010101110010100;
				12'h688: data <= 32'b00000000000000101010111001000001;
				12'h689: data <= 32'b00000000000000101011000011110001;
				12'h68A: data <= 32'b00000000000000101011001110100011;
				12'h68B: data <= 32'b00000000000000101011011001011000;
				12'h68C: data <= 32'b00000000000000101011100100001111;
				12'h68D: data <= 32'b00000000000000101011101111001010;
				12'h68E: data <= 32'b00000000000000101011111010000111;
				12'h68F: data <= 32'b00000000000000101100000101000111;
				12'h690: data <= 32'b00000000000000101100010000001010;
				12'h691: data <= 32'b00000000000000101100011011001111;
				12'h692: data <= 32'b00000000000000101100100110010111;
				12'h693: data <= 32'b00000000000000101100110001100010;
				12'h694: data <= 32'b00000000000000101100111100110000;
				12'h695: data <= 32'b00000000000000101101001000000001;
				12'h696: data <= 32'b00000000000000101101010011010100;
				12'h697: data <= 32'b00000000000000101101011110101010;
				12'h698: data <= 32'b00000000000000101101101010000011;
				12'h699: data <= 32'b00000000000000101101110101011111;
				12'h69A: data <= 32'b00000000000000101110000000111110;
				12'h69B: data <= 32'b00000000000000101110001100100000;
				12'h69C: data <= 32'b00000000000000101110011000000100;
				12'h69D: data <= 32'b00000000000000101110100011101100;
				12'h69E: data <= 32'b00000000000000101110101111010110;
				12'h69F: data <= 32'b00000000000000101110111011000100;
				12'h6A0: data <= 32'b00000000000000101111000110110100;
				12'h6A1: data <= 32'b00000000000000101111010010100111;
				12'h6A2: data <= 32'b00000000000000101111011110011101;
				12'h6A3: data <= 32'b00000000000000101111101010010110;
				12'h6A4: data <= 32'b00000000000000101111110110010010;
				12'h6A5: data <= 32'b00000000000000110000000010010001;
				12'h6A6: data <= 32'b00000000000000110000001110010011;
				12'h6A7: data <= 32'b00000000000000110000011010011001;
				12'h6A8: data <= 32'b00000000000000110000100110100001;
				12'h6A9: data <= 32'b00000000000000110000110010101100;
				12'h6AA: data <= 32'b00000000000000110000111110111010;
				12'h6AB: data <= 32'b00000000000000110001001011001011;
				12'h6AC: data <= 32'b00000000000000110001010111100000;
				12'h6AD: data <= 32'b00000000000000110001100011110111;
				12'h6AE: data <= 32'b00000000000000110001110000010001;
				12'h6AF: data <= 32'b00000000000000110001111100101111;
				12'h6B0: data <= 32'b00000000000000110010001001010000;
				12'h6B1: data <= 32'b00000000000000110010010101110100;
				12'h6B2: data <= 32'b00000000000000110010100010011011;
				12'h6B3: data <= 32'b00000000000000110010101111000101;
				12'h6B4: data <= 32'b00000000000000110010111011110010;
				12'h6B5: data <= 32'b00000000000000110011001000100011;
				12'h6B6: data <= 32'b00000000000000110011010101010111;
				12'h6B7: data <= 32'b00000000000000110011100010001110;
				12'h6B8: data <= 32'b00000000000000110011101111001000;
				12'h6B9: data <= 32'b00000000000000110011111100000101;
				12'h6BA: data <= 32'b00000000000000110100001001000110;
				12'h6BB: data <= 32'b00000000000000110100010110001010;
				12'h6BC: data <= 32'b00000000000000110100100011010001;
				12'h6BD: data <= 32'b00000000000000110100110000011011;
				12'h6BE: data <= 32'b00000000000000110100111101101001;
				12'h6BF: data <= 32'b00000000000000110101001010111010;
				12'h6C0: data <= 32'b00000000000000110101011000001111;
				12'h6C1: data <= 32'b00000000000000110101100101100110;
				12'h6C2: data <= 32'b00000000000000110101110011000001;
				12'h6C3: data <= 32'b00000000000000110110000000100000;
				12'h6C4: data <= 32'b00000000000000110110001110000010;
				12'h6C5: data <= 32'b00000000000000110110011011100111;
				12'h6C6: data <= 32'b00000000000000110110101001001111;
				12'h6C7: data <= 32'b00000000000000110110110110111011;
				12'h6C8: data <= 32'b00000000000000110111000100101011;
				12'h6C9: data <= 32'b00000000000000110111010010011110;
				12'h6CA: data <= 32'b00000000000000110111100000010100;
				12'h6CB: data <= 32'b00000000000000110111101110001110;
				12'h6CC: data <= 32'b00000000000000110111111100001011;
				12'h6CD: data <= 32'b00000000000000111000001010001100;
				12'h6CE: data <= 32'b00000000000000111000011000010000;
				12'h6CF: data <= 32'b00000000000000111000100110011000;
				12'h6D0: data <= 32'b00000000000000111000110100100100;
				12'h6D1: data <= 32'b00000000000000111001000010110010;
				12'h6D2: data <= 32'b00000000000000111001010001000101;
				12'h6D3: data <= 32'b00000000000000111001011111011011;
				12'h6D4: data <= 32'b00000000000000111001101101110101;
				12'h6D5: data <= 32'b00000000000000111001111100010010;
				12'h6D6: data <= 32'b00000000000000111010001010110011;
				12'h6D7: data <= 32'b00000000000000111010011001010111;
				12'h6D8: data <= 32'b00000000000000111010101000000000;
				12'h6D9: data <= 32'b00000000000000111010110110101011;
				12'h6DA: data <= 32'b00000000000000111011000101011011;
				12'h6DB: data <= 32'b00000000000000111011010100001110;
				12'h6DC: data <= 32'b00000000000000111011100011000101;
				12'h6DD: data <= 32'b00000000000000111011110010000000;
				12'h6DE: data <= 32'b00000000000000111100000000111110;
				12'h6DF: data <= 32'b00000000000000111100010000000000;
				12'h6E0: data <= 32'b00000000000000111100011111000110;
				12'h6E1: data <= 32'b00000000000000111100101110010000;
				12'h6E2: data <= 32'b00000000000000111100111101011101;
				12'h6E3: data <= 32'b00000000000000111101001100101110;
				12'h6E4: data <= 32'b00000000000000111101011100000011;
				12'h6E5: data <= 32'b00000000000000111101101011011100;
				12'h6E6: data <= 32'b00000000000000111101111010111001;
				12'h6E7: data <= 32'b00000000000000111110001010011010;
				12'h6E8: data <= 32'b00000000000000111110011001111110;
				12'h6E9: data <= 32'b00000000000000111110101001100111;
				12'h6EA: data <= 32'b00000000000000111110111001010011;
				12'h6EB: data <= 32'b00000000000000111111001001000100;
				12'h6EC: data <= 32'b00000000000000111111011000111000;
				12'h6ED: data <= 32'b00000000000000111111101000110000;
				12'h6EE: data <= 32'b00000000000000111111111000101100;
				12'h6EF: data <= 32'b00000000000001000000001000101100;
				12'h6F0: data <= 32'b00000000000001000000011000110001;
				12'h6F1: data <= 32'b00000000000001000000101000111001;
				12'h6F2: data <= 32'b00000000000001000000111001000101;
				12'h6F3: data <= 32'b00000000000001000001001001010101;
				12'h6F4: data <= 32'b00000000000001000001011001101010;
				12'h6F5: data <= 32'b00000000000001000001101010000010;
				12'h6F6: data <= 32'b00000000000001000001111010011111;
				12'h6F7: data <= 32'b00000000000001000010001010111111;
				12'h6F8: data <= 32'b00000000000001000010011011100100;
				12'h6F9: data <= 32'b00000000000001000010101100001101;
				12'h6FA: data <= 32'b00000000000001000010111100111010;
				12'h6FB: data <= 32'b00000000000001000011001101101100;
				12'h6FC: data <= 32'b00000000000001000011011110100001;
				12'h6FD: data <= 32'b00000000000001000011101111011011;
				12'h6FE: data <= 32'b00000000000001000100000000011001;
				12'h6FF: data <= 32'b00000000000001000100010001011011;
				12'h700: data <= 32'b00000000000001000100100010100010;
				12'h701: data <= 32'b00000000000001000100110011101100;
				12'h702: data <= 32'b00000000000001000101000100111011;
				12'h703: data <= 32'b00000000000001000101010110001111;
				12'h704: data <= 32'b00000000000001000101100111100111;
				12'h705: data <= 32'b00000000000001000101111001000011;
				12'h706: data <= 32'b00000000000001000110001010100011;
				12'h707: data <= 32'b00000000000001000110011100001000;
				12'h708: data <= 32'b00000000000001000110101101110001;
				12'h709: data <= 32'b00000000000001000110111111011111;
				12'h70A: data <= 32'b00000000000001000111010001010001;
				12'h70B: data <= 32'b00000000000001000111100011000111;
				12'h70C: data <= 32'b00000000000001000111110101000010;
				12'h70D: data <= 32'b00000000000001001000000111000010;
				12'h70E: data <= 32'b00000000000001001000011001000110;
				12'h70F: data <= 32'b00000000000001001000101011001111;
				12'h710: data <= 32'b00000000000001001000111101011100;
				12'h711: data <= 32'b00000000000001001001001111101101;
				12'h712: data <= 32'b00000000000001001001100010000100;
				12'h713: data <= 32'b00000000000001001001110100011110;
				12'h714: data <= 32'b00000000000001001010000110111110;
				12'h715: data <= 32'b00000000000001001010011001100010;
				12'h716: data <= 32'b00000000000001001010101100001011;
				12'h717: data <= 32'b00000000000001001010111110111000;
				12'h718: data <= 32'b00000000000001001011010001101010;
				12'h719: data <= 32'b00000000000001001011100100100001;
				12'h71A: data <= 32'b00000000000001001011110111011100;
				12'h71B: data <= 32'b00000000000001001100001010011100;
				12'h71C: data <= 32'b00000000000001001100011101100001;
				12'h71D: data <= 32'b00000000000001001100110000101011;
				12'h71E: data <= 32'b00000000000001001101000011111010;
				12'h71F: data <= 32'b00000000000001001101010111001101;
				12'h720: data <= 32'b00000000000001001101101010100101;
				12'h721: data <= 32'b00000000000001001101111110000011;
				12'h722: data <= 32'b00000000000001001110010001100100;
				12'h723: data <= 32'b00000000000001001110100101001011;
				12'h724: data <= 32'b00000000000001001110111000110111;
				12'h725: data <= 32'b00000000000001001111001100101000;
				12'h726: data <= 32'b00000000000001001111100000011101;
				12'h727: data <= 32'b00000000000001001111110100011000;
				12'h728: data <= 32'b00000000000001010000001000011000;
				12'h729: data <= 32'b00000000000001010000011100011100;
				12'h72A: data <= 32'b00000000000001010000110000100110;
				12'h72B: data <= 32'b00000000000001010001000100110100;
				12'h72C: data <= 32'b00000000000001010001011001001000;
				12'h72D: data <= 32'b00000000000001010001101101100001;
				12'h72E: data <= 32'b00000000000001010010000001111111;
				12'h72F: data <= 32'b00000000000001010010010110100010;
				12'h730: data <= 32'b00000000000001010010101011001010;
				12'h731: data <= 32'b00000000000001010010111111111000;
				12'h732: data <= 32'b00000000000001010011010100101010;
				12'h733: data <= 32'b00000000000001010011101001100010;
				12'h734: data <= 32'b00000000000001010011111110011111;
				12'h735: data <= 32'b00000000000001010100010011100001;
				12'h736: data <= 32'b00000000000001010100101000101001;
				12'h737: data <= 32'b00000000000001010100111101110110;
				12'h738: data <= 32'b00000000000001010101010011001000;
				12'h739: data <= 32'b00000000000001010101101000011111;
				12'h73A: data <= 32'b00000000000001010101111101111100;
				12'h73B: data <= 32'b00000000000001010110010011011110;
				12'h73C: data <= 32'b00000000000001010110101001000110;
				12'h73D: data <= 32'b00000000000001010110111110110011;
				12'h73E: data <= 32'b00000000000001010111010100100101;
				12'h73F: data <= 32'b00000000000001010111101010011101;
				12'h740: data <= 32'b00000000000001011000000000011010;
				12'h741: data <= 32'b00000000000001011000010110011101;
				12'h742: data <= 32'b00000000000001011000101100100110;
				12'h743: data <= 32'b00000000000001011001000010110100;
				12'h744: data <= 32'b00000000000001011001011001000111;
				12'h745: data <= 32'b00000000000001011001101111100000;
				12'h746: data <= 32'b00000000000001011010000101111111;
				12'h747: data <= 32'b00000000000001011010011100100011;
				12'h748: data <= 32'b00000000000001011010110011001101;
				12'h749: data <= 32'b00000000000001011011001001111101;
				12'h74A: data <= 32'b00000000000001011011100000110010;
				12'h74B: data <= 32'b00000000000001011011110111101101;
				12'h74C: data <= 32'b00000000000001011100001110101110;
				12'h74D: data <= 32'b00000000000001011100100101110100;
				12'h74E: data <= 32'b00000000000001011100111101000001;
				12'h74F: data <= 32'b00000000000001011101010100010011;
				12'h750: data <= 32'b00000000000001011101101011101011;
				12'h751: data <= 32'b00000000000001011110000011001001;
				12'h752: data <= 32'b00000000000001011110011010101101;
				12'h753: data <= 32'b00000000000001011110110010010110;
				12'h754: data <= 32'b00000000000001011111001010000110;
				12'h755: data <= 32'b00000000000001011111100001111011;
				12'h756: data <= 32'b00000000000001011111111001110111;
				12'h757: data <= 32'b00000000000001100000010001111000;
				12'h758: data <= 32'b00000000000001100000101010000000;
				12'h759: data <= 32'b00000000000001100001000010001101;
				12'h75A: data <= 32'b00000000000001100001011010100001;
				12'h75B: data <= 32'b00000000000001100001110010111010;
				12'h75C: data <= 32'b00000000000001100010001011011010;
				12'h75D: data <= 32'b00000000000001100010100100000000;
				12'h75E: data <= 32'b00000000000001100010111100101100;
				12'h75F: data <= 32'b00000000000001100011010101011111;
				12'h760: data <= 32'b00000000000001100011101110010111;
				12'h761: data <= 32'b00000000000001100100000111010110;
				12'h762: data <= 32'b00000000000001100100100000011011;
				12'h763: data <= 32'b00000000000001100100111001100110;
				12'h764: data <= 32'b00000000000001100101010010110111;
				12'h765: data <= 32'b00000000000001100101101100001111;
				12'h766: data <= 32'b00000000000001100110000101101110;
				12'h767: data <= 32'b00000000000001100110011111010010;
				12'h768: data <= 32'b00000000000001100110111000111101;
				12'h769: data <= 32'b00000000000001100111010010101111;
				12'h76A: data <= 32'b00000000000001100111101100100111;
				12'h76B: data <= 32'b00000000000001101000000110100101;
				12'h76C: data <= 32'b00000000000001101000100000101010;
				12'h76D: data <= 32'b00000000000001101000111010110101;
				12'h76E: data <= 32'b00000000000001101001010101000111;
				12'h76F: data <= 32'b00000000000001101001101111100000;
				12'h770: data <= 32'b00000000000001101010001001111111;
				12'h771: data <= 32'b00000000000001101010100100100101;
				12'h772: data <= 32'b00000000000001101010111111010001;
				12'h773: data <= 32'b00000000000001101011011010000101;
				12'h774: data <= 32'b00000000000001101011110100111111;
				12'h775: data <= 32'b00000000000001101100001111111111;
				12'h776: data <= 32'b00000000000001101100101011000111;
				12'h777: data <= 32'b00000000000001101101000110010101;
				12'h778: data <= 32'b00000000000001101101100001101010;
				12'h779: data <= 32'b00000000000001101101111101000110;
				12'h77A: data <= 32'b00000000000001101110011000101000;
				12'h77B: data <= 32'b00000000000001101110110100010010;
				12'h77C: data <= 32'b00000000000001101111010000000010;
				12'h77D: data <= 32'b00000000000001101111101011111010;
				12'h77E: data <= 32'b00000000000001110000000111111000;
				12'h77F: data <= 32'b00000000000001110000100011111110;
				12'h780: data <= 32'b00000000000001110001000000001010;
				12'h781: data <= 32'b00000000000001110001011100011110;
				12'h782: data <= 32'b00000000000001110001111000111001;
				12'h783: data <= 32'b00000000000001110010010101011010;
				12'h784: data <= 32'b00000000000001110010110010000011;
				12'h785: data <= 32'b00000000000001110011001110110011;
				12'h786: data <= 32'b00000000000001110011101011101011;
				12'h787: data <= 32'b00000000000001110100001000101001;
				12'h788: data <= 32'b00000000000001110100100101101111;
				12'h789: data <= 32'b00000000000001110101000010111100;
				12'h78A: data <= 32'b00000000000001110101100000010001;
				12'h78B: data <= 32'b00000000000001110101111101101100;
				12'h78C: data <= 32'b00000000000001110110011011001111;
				12'h78D: data <= 32'b00000000000001110110111000111010;
				12'h78E: data <= 32'b00000000000001110111010110101100;
				12'h78F: data <= 32'b00000000000001110111110100100101;
				12'h790: data <= 32'b00000000000001111000010010100110;
				12'h791: data <= 32'b00000000000001111000110000101111;
				12'h792: data <= 32'b00000000000001111001001110111111;
				12'h793: data <= 32'b00000000000001111001101101010110;
				12'h794: data <= 32'b00000000000001111010001011110101;
				12'h795: data <= 32'b00000000000001111010101010011100;
				12'h796: data <= 32'b00000000000001111011001001001010;
				12'h797: data <= 32'b00000000000001111011101000000001;
				12'h798: data <= 32'b00000000000001111100000110111111;
				12'h799: data <= 32'b00000000000001111100100110000100;
				12'h79A: data <= 32'b00000000000001111101000101010010;
				12'h79B: data <= 32'b00000000000001111101100100100111;
				12'h79C: data <= 32'b00000000000001111110000100000100;
				12'h79D: data <= 32'b00000000000001111110100011101001;
				12'h79E: data <= 32'b00000000000001111111000011010110;
				12'h79F: data <= 32'b00000000000001111111100011001011;
				12'h7A0: data <= 32'b00000000000010000000000011000111;
				12'h7A1: data <= 32'b00000000000010000000100011001100;
				12'h7A2: data <= 32'b00000000000010000001000011011001;
				12'h7A3: data <= 32'b00000000000010000001100011101110;
				12'h7A4: data <= 32'b00000000000010000010000100001011;
				12'h7A5: data <= 32'b00000000000010000010100100110000;
				12'h7A6: data <= 32'b00000000000010000011000101011101;
				12'h7A7: data <= 32'b00000000000010000011100110010011;
				12'h7A8: data <= 32'b00000000000010000100000111010000;
				12'h7A9: data <= 32'b00000000000010000100101000010110;
				12'h7AA: data <= 32'b00000000000010000101001001100101;
				12'h7AB: data <= 32'b00000000000010000101101010111011;
				12'h7AC: data <= 32'b00000000000010000110001100011010;
				12'h7AD: data <= 32'b00000000000010000110101110000001;
				12'h7AE: data <= 32'b00000000000010000111001111110001;
				12'h7AF: data <= 32'b00000000000010000111110001101001;
				12'h7B0: data <= 32'b00000000000010001000010011101010;
				12'h7B1: data <= 32'b00000000000010001000110101110011;
				12'h7B2: data <= 32'b00000000000010001001011000000101;
				12'h7B3: data <= 32'b00000000000010001001111010011111;
				12'h7B4: data <= 32'b00000000000010001010011101000010;
				12'h7B5: data <= 32'b00000000000010001010111111101110;
				12'h7B6: data <= 32'b00000000000010001011100010100010;
				12'h7B7: data <= 32'b00000000000010001100000101011111;
				12'h7B8: data <= 32'b00000000000010001100101000100101;
				12'h7B9: data <= 32'b00000000000010001101001011110011;
				12'h7BA: data <= 32'b00000000000010001101101111001011;
				12'h7BB: data <= 32'b00000000000010001110010010101011;
				12'h7BC: data <= 32'b00000000000010001110110110010100;
				12'h7BD: data <= 32'b00000000000010001111011010000110;
				12'h7BE: data <= 32'b00000000000010001111111110000001;
				12'h7BF: data <= 32'b00000000000010010000100010000101;
				12'h7C0: data <= 32'b00000000000010010001000110010010;
				12'h7C1: data <= 32'b00000000000010010001101010101000;
				12'h7C2: data <= 32'b00000000000010010010001111000111;
				12'h7C3: data <= 32'b00000000000010010010110011110000;
				12'h7C4: data <= 32'b00000000000010010011011000100001;
				12'h7C5: data <= 32'b00000000000010010011111101011100;
				12'h7C6: data <= 32'b00000000000010010100100010100000;
				12'h7C7: data <= 32'b00000000000010010101000111101101;
				12'h7C8: data <= 32'b00000000000010010101101101000100;
				12'h7C9: data <= 32'b00000000000010010110010010100100;
				12'h7CA: data <= 32'b00000000000010010110111000001101;
				12'h7CB: data <= 32'b00000000000010010111011110000000;
				12'h7CC: data <= 32'b00000000000010011000000011111100;
				12'h7CD: data <= 32'b00000000000010011000101010000010;
				12'h7CE: data <= 32'b00000000000010011001010000010001;
				12'h7CF: data <= 32'b00000000000010011001110110101010;
				12'h7D0: data <= 32'b00000000000010011010011101001101;
				12'h7D1: data <= 32'b00000000000010011011000011111001;
				12'h7D2: data <= 32'b00000000000010011011101010101111;
				12'h7D3: data <= 32'b00000000000010011100010001101110;
				12'h7D4: data <= 32'b00000000000010011100111000110111;
				12'h7D5: data <= 32'b00000000000010011101100000001011;
				12'h7D6: data <= 32'b00000000000010011110000111100111;
				12'h7D7: data <= 32'b00000000000010011110101111001110;
				12'h7D8: data <= 32'b00000000000010011111010110111111;
				12'h7D9: data <= 32'b00000000000010011111111110111010;
				12'h7DA: data <= 32'b00000000000010100000100110111111;
				12'h7DB: data <= 32'b00000000000010100001001111001101;
				12'h7DC: data <= 32'b00000000000010100001110111100110;
				12'h7DD: data <= 32'b00000000000010100010100000001001;
				12'h7DE: data <= 32'b00000000000010100011001000110110;
				12'h7DF: data <= 32'b00000000000010100011110001101110;
				12'h7E0: data <= 32'b00000000000010100100011010101111;
				12'h7E1: data <= 32'b00000000000010100101000011111011;
				12'h7E2: data <= 32'b00000000000010100101101101010001;
				12'h7E3: data <= 32'b00000000000010100110010110110010;
				12'h7E4: data <= 32'b00000000000010100111000000011101;
				12'h7E5: data <= 32'b00000000000010100111101010010010;
				12'h7E6: data <= 32'b00000000000010101000010100010010;
				12'h7E7: data <= 32'b00000000000010101000111110011100;
				12'h7E8: data <= 32'b00000000000010101001101000110001;
				12'h7E9: data <= 32'b00000000000010101010010011010000;
				12'h7EA: data <= 32'b00000000000010101010111101111011;
				12'h7EB: data <= 32'b00000000000010101011101000101111;
				12'h7EC: data <= 32'b00000000000010101100010011101111;
				12'h7ED: data <= 32'b00000000000010101100111110111001;
				12'h7EE: data <= 32'b00000000000010101101101010001110;
				12'h7EF: data <= 32'b00000000000010101110010101101110;
				12'h7F0: data <= 32'b00000000000010101111000001011001;
				12'h7F1: data <= 32'b00000000000010101111101101001111;
				12'h7F2: data <= 32'b00000000000010110000011001010000;
				12'h7F3: data <= 32'b00000000000010110001000101011100;
				12'h7F4: data <= 32'b00000000000010110001110001110011;
				12'h7F5: data <= 32'b00000000000010110010011110010101;
				12'h7F6: data <= 32'b00000000000010110011001011000010;
				12'h7F7: data <= 32'b00000000000010110011110111111010;
				12'h7F8: data <= 32'b00000000000010110100100100111110;
				12'h7F9: data <= 32'b00000000000010110101010010001101;
				12'h7FA: data <= 32'b00000000000010110101111111100111;
				12'h7FB: data <= 32'b00000000000010110110101101001101;
				12'h7FC: data <= 32'b00000000000010110111011010111110;
				12'h7FD: data <= 32'b00000000000010111000001000111010;
				12'h7FE: data <= 32'b00000000000010111000110111000010;
				12'h7FF: data <= 32'b00000000000010111001100101010110;
				12'h800: data <= 32'b00000000000010111010010011110101;
				12'h801: data <= 32'b00000000000010111011000010100000;
				12'h802: data <= 32'b00000000000010111011110001010110;
				12'h803: data <= 32'b00000000000010111100100000011000;
				12'h804: data <= 32'b00000000000010111101001111100110;
				12'h805: data <= 32'b00000000000010111101111111000000;
				12'h806: data <= 32'b00000000000010111110101110100110;
				12'h807: data <= 32'b00000000000010111111011110010111;
				12'h808: data <= 32'b00000000000011000000001110010101;
				12'h809: data <= 32'b00000000000011000000111110011111;
				12'h80A: data <= 32'b00000000000011000001101110110100;
				12'h80B: data <= 32'b00000000000011000010011111010110;
				12'h80C: data <= 32'b00000000000011000011010000000100;
				12'h80D: data <= 32'b00000000000011000100000000111110;
				12'h80E: data <= 32'b00000000000011000100110010000100;
				12'h80F: data <= 32'b00000000000011000101100011010111;
				12'h810: data <= 32'b00000000000011000110010100110110;
				12'h811: data <= 32'b00000000000011000111000110100010;
				12'h812: data <= 32'b00000000000011000111111000011001;
				12'h813: data <= 32'b00000000000011001000101010011110;
				12'h814: data <= 32'b00000000000011001001011100101111;
				12'h815: data <= 32'b00000000000011001010001111001100;
				12'h816: data <= 32'b00000000000011001011000001110110;
				12'h817: data <= 32'b00000000000011001011110100101101;
				12'h818: data <= 32'b00000000000011001100100111110001;
				12'h819: data <= 32'b00000000000011001101011011000001;
				12'h81A: data <= 32'b00000000000011001110001110011110;
				12'h81B: data <= 32'b00000000000011001111000010001000;
				12'h81C: data <= 32'b00000000000011001111110101111111;
				12'h81D: data <= 32'b00000000000011010000101010000011;
				12'h81E: data <= 32'b00000000000011010001011110010100;
				12'h81F: data <= 32'b00000000000011010010010010110010;
				12'h820: data <= 32'b00000000000011010011000111011110;
				12'h821: data <= 32'b00000000000011010011111100010110;
				12'h822: data <= 32'b00000000000011010100110001011100;
				12'h823: data <= 32'b00000000000011010101100110101111;
				12'h824: data <= 32'b00000000000011010110011100001111;
				12'h825: data <= 32'b00000000000011010111010001111101;
				12'h826: data <= 32'b00000000000011011000000111111000;
				12'h827: data <= 32'b00000000000011011000111110000001;
				12'h828: data <= 32'b00000000000011011001110100010111;
				12'h829: data <= 32'b00000000000011011010101010111011;
				12'h82A: data <= 32'b00000000000011011011100001101101;
				12'h82B: data <= 32'b00000000000011011100011000101100;
				12'h82C: data <= 32'b00000000000011011101001111111001;
				12'h82D: data <= 32'b00000000000011011110000111010100;
				12'h82E: data <= 32'b00000000000011011110111110111101;
				12'h82F: data <= 32'b00000000000011011111110110110100;
				12'h830: data <= 32'b00000000000011100000101110111000;
				12'h831: data <= 32'b00000000000011100001100111001011;
				12'h832: data <= 32'b00000000000011100010011111101100;
				12'h833: data <= 32'b00000000000011100011011000011011;
				12'h834: data <= 32'b00000000000011100100010001011000;
				12'h835: data <= 32'b00000000000011100101001010100100;
				12'h836: data <= 32'b00000000000011100110000011111101;
				12'h837: data <= 32'b00000000000011100110111101100110;
				12'h838: data <= 32'b00000000000011100111110111011100;
				12'h839: data <= 32'b00000000000011101000110001100001;
				12'h83A: data <= 32'b00000000000011101001101011110101;
				12'h83B: data <= 32'b00000000000011101010100110010111;
				12'h83C: data <= 32'b00000000000011101011100001001000;
				12'h83D: data <= 32'b00000000000011101100011100001000;
				12'h83E: data <= 32'b00000000000011101101010111010110;
				12'h83F: data <= 32'b00000000000011101110010010110100;
				12'h840: data <= 32'b00000000000011101111001110100000;
				12'h841: data <= 32'b00000000000011110000001010011011;
				12'h842: data <= 32'b00000000000011110001000110100101;
				12'h843: data <= 32'b00000000000011110010000010111110;
				12'h844: data <= 32'b00000000000011110010111111100110;
				12'h845: data <= 32'b00000000000011110011111100011110;
				12'h846: data <= 32'b00000000000011110100111001100101;
				12'h847: data <= 32'b00000000000011110101110110111011;
				12'h848: data <= 32'b00000000000011110110110100100000;
				12'h849: data <= 32'b00000000000011110111110010010101;
				12'h84A: data <= 32'b00000000000011111000110000011001;
				12'h84B: data <= 32'b00000000000011111001101110101101;
				12'h84C: data <= 32'b00000000000011111010101101010001;
				12'h84D: data <= 32'b00000000000011111011101100000100;
				12'h84E: data <= 32'b00000000000011111100101011000111;
				12'h84F: data <= 32'b00000000000011111101101010011001;
				12'h850: data <= 32'b00000000000011111110101001111100;
				12'h851: data <= 32'b00000000000011111111101001101110;
				12'h852: data <= 32'b00000000000100000000101001110001;
				12'h853: data <= 32'b00000000000100000001101010000011;
				12'h854: data <= 32'b00000000000100000010101010100110;
				12'h855: data <= 32'b00000000000100000011101011011001;
				12'h856: data <= 32'b00000000000100000100101100011100;
				12'h857: data <= 32'b00000000000100000101101101101111;
				12'h858: data <= 32'b00000000000100000110101111010011;
				12'h859: data <= 32'b00000000000100000111110001000111;
				12'h85A: data <= 32'b00000000000100001000110011001011;
				12'h85B: data <= 32'b00000000000100001001110101100000;
				12'h85C: data <= 32'b00000000000100001010111000000110;
				12'h85D: data <= 32'b00000000000100001011111010111100;
				12'h85E: data <= 32'b00000000000100001100111110000011;
				12'h85F: data <= 32'b00000000000100001110000001011011;
				12'h860: data <= 32'b00000000000100001111000101000100;
				12'h861: data <= 32'b00000000000100010000001000111110;
				12'h862: data <= 32'b00000000000100010001001101001001;
				12'h863: data <= 32'b00000000000100010010010001100101;
				12'h864: data <= 32'b00000000000100010011010110010010;
				12'h865: data <= 32'b00000000000100010100011011010000;
				12'h866: data <= 32'b00000000000100010101100000011111;
				12'h867: data <= 32'b00000000000100010110100110000000;
				12'h868: data <= 32'b00000000000100010111101011110010;
				12'h869: data <= 32'b00000000000100011000110001110110;
				12'h86A: data <= 32'b00000000000100011001111000001011;
				12'h86B: data <= 32'b00000000000100011010111110110010;
				12'h86C: data <= 32'b00000000000100011100000101101011;
				12'h86D: data <= 32'b00000000000100011101001100110101;
				12'h86E: data <= 32'b00000000000100011110010100010001;
				12'h86F: data <= 32'b00000000000100011111011011111111;
				12'h870: data <= 32'b00000000000100100000100011111111;
				12'h871: data <= 32'b00000000000100100001101100010001;
				12'h872: data <= 32'b00000000000100100010110100110101;
				12'h873: data <= 32'b00000000000100100011111101101011;
				12'h874: data <= 32'b00000000000100100101000110110100;
				12'h875: data <= 32'b00000000000100100110010000001111;
				12'h876: data <= 32'b00000000000100100111011001111100;
				12'h877: data <= 32'b00000000000100101000100011111100;
				12'h878: data <= 32'b00000000000100101001101110001110;
				12'h879: data <= 32'b00000000000100101010111000110011;
				12'h87A: data <= 32'b00000000000100101100000011101011;
				12'h87B: data <= 32'b00000000000100101101001110110101;
				12'h87C: data <= 32'b00000000000100101110011010010010;
				12'h87D: data <= 32'b00000000000100101111100110000010;
				12'h87E: data <= 32'b00000000000100110000110010000101;
				12'h87F: data <= 32'b00000000000100110001111110011011;
				12'h880: data <= 32'b00000000000100110011001011000100;
				12'h881: data <= 32'b00000000000100110100011000000001;
				12'h882: data <= 32'b00000000000100110101100101010000;
				12'h883: data <= 32'b00000000000100110110110010110011;
				12'h884: data <= 32'b00000000000100111000000000101010;
				12'h885: data <= 32'b00000000000100111001001110110100;
				12'h886: data <= 32'b00000000000100111010011101010001;
				12'h887: data <= 32'b00000000000100111011101100000010;
				12'h888: data <= 32'b00000000000100111100111011000111;
				12'h889: data <= 32'b00000000000100111110001010100000;
				12'h88A: data <= 32'b00000000000100111111011010001101;
				12'h88B: data <= 32'b00000000000101000000101010001101;
				12'h88C: data <= 32'b00000000000101000001111010100010;
				12'h88D: data <= 32'b00000000000101000011001011001010;
				12'h88E: data <= 32'b00000000000101000100011100000111;
				12'h88F: data <= 32'b00000000000101000101101101011000;
				12'h890: data <= 32'b00000000000101000110111110111110;
				12'h891: data <= 32'b00000000000101001000010000111000;
				12'h892: data <= 32'b00000000000101001001100011000110;
				12'h893: data <= 32'b00000000000101001010110101101010;
				12'h894: data <= 32'b00000000000101001100001000100001;
				12'h895: data <= 32'b00000000000101001101011011101110;
				12'h896: data <= 32'b00000000000101001110101111001111;
				12'h897: data <= 32'b00000000000101010000000011000110;
				12'h898: data <= 32'b00000000000101010001010111010001;
				12'h899: data <= 32'b00000000000101010010101011110001;
				12'h89A: data <= 32'b00000000000101010100000000100111;
				12'h89B: data <= 32'b00000000000101010101010101110010;
				12'h89C: data <= 32'b00000000000101010110101011010010;
				12'h89D: data <= 32'b00000000000101011000000001000111;
				12'h89E: data <= 32'b00000000000101011001010111010010;
				12'h89F: data <= 32'b00000000000101011010101101110011;
				12'h8A0: data <= 32'b00000000000101011100000100101001;
				12'h8A1: data <= 32'b00000000000101011101011011110101;
				12'h8A2: data <= 32'b00000000000101011110110011010111;
				12'h8A3: data <= 32'b00000000000101100000001011001111;
				12'h8A4: data <= 32'b00000000000101100001100011011101;
				12'h8A5: data <= 32'b00000000000101100010111100000001;
				12'h8A6: data <= 32'b00000000000101100100010100111011;
				12'h8A7: data <= 32'b00000000000101100101101110001011;
				12'h8A8: data <= 32'b00000000000101100111000111110010;
				12'h8A9: data <= 32'b00000000000101101000100001101111;
				12'h8AA: data <= 32'b00000000000101101001111100000011;
				12'h8AB: data <= 32'b00000000000101101011010110101101;
				12'h8AC: data <= 32'b00000000000101101100110001101110;
				12'h8AD: data <= 32'b00000000000101101110001101000110;
				12'h8AE: data <= 32'b00000000000101101111101000110101;
				12'h8AF: data <= 32'b00000000000101110001000100111010;
				12'h8B0: data <= 32'b00000000000101110010100001010111;
				12'h8B1: data <= 32'b00000000000101110011111110001011;
				12'h8B2: data <= 32'b00000000000101110101011011010110;
				12'h8B3: data <= 32'b00000000000101110110111000111001;
				12'h8B4: data <= 32'b00000000000101111000010110110011;
				12'h8B5: data <= 32'b00000000000101111001110101000100;
				12'h8B6: data <= 32'b00000000000101111011010011101101;
				12'h8B7: data <= 32'b00000000000101111100110010101110;
				12'h8B8: data <= 32'b00000000000101111110010010000111;
				12'h8B9: data <= 32'b00000000000101111111110001110111;
				12'h8BA: data <= 32'b00000000000110000001010010000000;
				12'h8BB: data <= 32'b00000000000110000010110010100000;
				12'h8BC: data <= 32'b00000000000110000100010011011001;
				12'h8BD: data <= 32'b00000000000110000101110100101010;
				12'h8BE: data <= 32'b00000000000110000111010110010011;
				12'h8BF: data <= 32'b00000000000110001000111000010101;
				12'h8C0: data <= 32'b00000000000110001010011010110000;
				12'h8C1: data <= 32'b00000000000110001011111101100011;
				12'h8C2: data <= 32'b00000000000110001101100000101110;
				12'h8C3: data <= 32'b00000000000110001111000100010011;
				12'h8C4: data <= 32'b00000000000110010000101000010001;
				12'h8C5: data <= 32'b00000000000110010010001100100111;
				12'h8C6: data <= 32'b00000000000110010011110001010111;
				12'h8C7: data <= 32'b00000000000110010101010110100000;
				12'h8C8: data <= 32'b00000000000110010110111100000010;
				12'h8C9: data <= 32'b00000000000110011000100001111110;
				12'h8CA: data <= 32'b00000000000110011010001000010011;
				12'h8CB: data <= 32'b00000000000110011011101111000010;
				12'h8CC: data <= 32'b00000000000110011101010110001011;
				12'h8CD: data <= 32'b00000000000110011110111101101101;
				12'h8CE: data <= 32'b00000000000110100000100101101010;
				12'h8CF: data <= 32'b00000000000110100010001110000000;
				12'h8D0: data <= 32'b00000000000110100011110110110001;
				12'h8D1: data <= 32'b00000000000110100101011111111100;
				12'h8D2: data <= 32'b00000000000110100111001001100001;
				12'h8D3: data <= 32'b00000000000110101000110011100000;
				12'h8D4: data <= 32'b00000000000110101010011101111011;
				12'h8D5: data <= 32'b00000000000110101100001000101111;
				12'h8D6: data <= 32'b00000000000110101101110011111111;
				12'h8D7: data <= 32'b00000000000110101111011111101001;
				12'h8D8: data <= 32'b00000000000110110001001011101111;
				12'h8D9: data <= 32'b00000000000110110010111000001111;
				12'h8DA: data <= 32'b00000000000110110100100101001011;
				12'h8DB: data <= 32'b00000000000110110110010010100010;
				12'h8DC: data <= 32'b00000000000110111000000000010100;
				12'h8DD: data <= 32'b00000000000110111001101110100010;
				12'h8DE: data <= 32'b00000000000110111011011101001100;
				12'h8DF: data <= 32'b00000000000110111101001100010001;
				12'h8E0: data <= 32'b00000000000110111110111011110010;
				12'h8E1: data <= 32'b00000000000111000000101011101111;
				12'h8E2: data <= 32'b00000000000111000010011100001000;
				12'h8E3: data <= 32'b00000000000111000100001100111101;
				12'h8E4: data <= 32'b00000000000111000101111110001110;
				12'h8E5: data <= 32'b00000000000111000111101111111100;
				12'h8E6: data <= 32'b00000000000111001001100010000110;
				12'h8E7: data <= 32'b00000000000111001011010100101101;
				12'h8E8: data <= 32'b00000000000111001101000111110001;
				12'h8E9: data <= 32'b00000000000111001110111011010001;
				12'h8EA: data <= 32'b00000000000111010000101111001110;
				12'h8EB: data <= 32'b00000000000111010010100011101001;
				12'h8EC: data <= 32'b00000000000111010100011000100000;
				12'h8ED: data <= 32'b00000000000111010110001101110101;
				12'h8EE: data <= 32'b00000000000111011000000011100111;
				12'h8EF: data <= 32'b00000000000111011001111001110111;
				12'h8F0: data <= 32'b00000000000111011011110000100100;
				12'h8F1: data <= 32'b00000000000111011101100111101111;
				12'h8F2: data <= 32'b00000000000111011111011111011000;
				12'h8F3: data <= 32'b00000000000111100001010111011111;
				12'h8F4: data <= 32'b00000000000111100011010000000100;
				12'h8F5: data <= 32'b00000000000111100101001001000111;
				12'h8F6: data <= 32'b00000000000111100111000010101000;
				12'h8F7: data <= 32'b00000000000111101000111100101000;
				12'h8F8: data <= 32'b00000000000111101010110111000111;
				12'h8F9: data <= 32'b00000000000111101100110010000100;
				12'h8FA: data <= 32'b00000000000111101110101101100000;
				12'h8FB: data <= 32'b00000000000111110000101001011011;
				12'h8FC: data <= 32'b00000000000111110010100101110101;
				12'h8FD: data <= 32'b00000000000111110100100010101110;
				12'h8FE: data <= 32'b00000000000111110110100000000110;
				12'h8FF: data <= 32'b00000000000111111000011101111110;
				12'h900: data <= 32'b00000000000111111010011100010101;
				12'h901: data <= 32'b00000000000111111100011011001100;
				12'h902: data <= 32'b00000000000111111110011010100011;
				12'h903: data <= 32'b00000000001000000000011010011001;
				12'h904: data <= 32'b00000000001000000010011010110000;
				12'h905: data <= 32'b00000000001000000100011011100111;
				12'h906: data <= 32'b00000000001000000110011100111110;
				12'h907: data <= 32'b00000000001000001000011110110101;
				12'h908: data <= 32'b00000000001000001010100001001101;
				12'h909: data <= 32'b00000000001000001100100100000110;
				12'h90A: data <= 32'b00000000001000001110100111011111;
				12'h90B: data <= 32'b00000000001000010000101011011010;
				12'h90C: data <= 32'b00000000001000010010101111110101;
				12'h90D: data <= 32'b00000000001000010100110100110010;
				12'h90E: data <= 32'b00000000001000010110111010001111;
				12'h90F: data <= 32'b00000000001000011001000000001111;
				12'h910: data <= 32'b00000000001000011011000110110000;
				12'h911: data <= 32'b00000000001000011101001101110010;
				12'h912: data <= 32'b00000000001000011111010101010111;
				12'h913: data <= 32'b00000000001000100001011101011101;
				12'h914: data <= 32'b00000000001000100011100110000101;
				12'h915: data <= 32'b00000000001000100101101111010000;
				12'h916: data <= 32'b00000000001000100111111000111101;
				12'h917: data <= 32'b00000000001000101010000011001101;
				12'h918: data <= 32'b00000000001000101100001101111111;
				12'h919: data <= 32'b00000000001000101110011001010100;
				12'h91A: data <= 32'b00000000001000110000100101001011;
				12'h91B: data <= 32'b00000000001000110010110001100110;
				12'h91C: data <= 32'b00000000001000110100111110100100;
				12'h91D: data <= 32'b00000000001000110111001100000110;
				12'h91E: data <= 32'b00000000001000111001011010001010;
				12'h91F: data <= 32'b00000000001000111011101000110011;
				12'h920: data <= 32'b00000000001000111101110111111111;
				12'h921: data <= 32'b00000000001001000000000111101111;
				12'h922: data <= 32'b00000000001001000010011000000011;
				12'h923: data <= 32'b00000000001001000100101000111011;
				12'h924: data <= 32'b00000000001001000110111010010111;
				12'h925: data <= 32'b00000000001001001001001100011000;
				12'h926: data <= 32'b00000000001001001011011110111101;
				12'h927: data <= 32'b00000000001001001101110010001000;
				12'h928: data <= 32'b00000000001001010000000101110111;
				12'h929: data <= 32'b00000000001001010010011010001011;
				12'h92A: data <= 32'b00000000001001010100101111000100;
				12'h92B: data <= 32'b00000000001001010111000100100010;
				12'h92C: data <= 32'b00000000001001011001011010100110;
				12'h92D: data <= 32'b00000000001001011011110001001111;
				12'h92E: data <= 32'b00000000001001011110001000011111;
				12'h92F: data <= 32'b00000000001001100000100000010100;
				12'h930: data <= 32'b00000000001001100010111000101111;
				12'h931: data <= 32'b00000000001001100101010001110000;
				12'h932: data <= 32'b00000000001001100111101011011000;
				12'h933: data <= 32'b00000000001001101010000101100110;
				12'h934: data <= 32'b00000000001001101100100000011011;
				12'h935: data <= 32'b00000000001001101110111011110110;
				12'h936: data <= 32'b00000000001001110001010111111001;
				12'h937: data <= 32'b00000000001001110011110100100010;
				12'h938: data <= 32'b00000000001001110110010001110011;
				12'h939: data <= 32'b00000000001001111000101111101011;
				12'h93A: data <= 32'b00000000001001111011001110001011;
				12'h93B: data <= 32'b00000000001001111101101101010010;
				12'h93C: data <= 32'b00000000001010000000001101000010;
				12'h93D: data <= 32'b00000000001010000010101101011001;
				12'h93E: data <= 32'b00000000001010000101001110011000;
				12'h93F: data <= 32'b00000000001010000111110000000000;
				12'h940: data <= 32'b00000000001010001010010010010000;
				12'h941: data <= 32'b00000000001010001100110101001001;
				12'h942: data <= 32'b00000000001010001111011000101011;
				12'h943: data <= 32'b00000000001010010001111100110110;
				12'h944: data <= 32'b00000000001010010100100001101001;
				12'h945: data <= 32'b00000000001010010111000111000111;
				12'h946: data <= 32'b00000000001010011001101101001101;
				12'h947: data <= 32'b00000000001010011100010011111101;
				12'h948: data <= 32'b00000000001010011110111011010111;
				12'h949: data <= 32'b00000000001010100001100011011011;
				12'h94A: data <= 32'b00000000001010100100001100001001;
				12'h94B: data <= 32'b00000000001010100110110101100001;
				12'h94C: data <= 32'b00000000001010101001011111100100;
				12'h94D: data <= 32'b00000000001010101100001010010001;
				12'h94E: data <= 32'b00000000001010101110110101101001;
				12'h94F: data <= 32'b00000000001010110001100001101100;
				12'h950: data <= 32'b00000000001010110100001110011010;
				12'h951: data <= 32'b00000000001010110110111011110011;
				12'h952: data <= 32'b00000000001010111001101001111000;
				12'h953: data <= 32'b00000000001010111100011000101000;
				12'h954: data <= 32'b00000000001010111111001000000100;
				12'h955: data <= 32'b00000000001011000001111000001100;
				12'h956: data <= 32'b00000000001011000100101001000000;
				12'h957: data <= 32'b00000000001011000111011010100001;
				12'h958: data <= 32'b00000000001011001010001100101110;
				12'h959: data <= 32'b00000000001011001100111111100111;
				12'h95A: data <= 32'b00000000001011001111110011001101;
				12'h95B: data <= 32'b00000000001011010010100111100001;
				12'h95C: data <= 32'b00000000001011010101011100100001;
				12'h95D: data <= 32'b00000000001011011000010010001111;
				12'h95E: data <= 32'b00000000001011011011001000101010;
				12'h95F: data <= 32'b00000000001011011101111111110011;
				12'h960: data <= 32'b00000000001011100000110111101010;
				12'h961: data <= 32'b00000000001011100011110000001111;
				12'h962: data <= 32'b00000000001011100110101001100011;
				12'h963: data <= 32'b00000000001011101001100011100100;
				12'h964: data <= 32'b00000000001011101100011110010100;
				12'h965: data <= 32'b00000000001011101111011001110011;
				12'h966: data <= 32'b00000000001011110010010110000001;
				12'h967: data <= 32'b00000000001011110101010010111111;
				12'h968: data <= 32'b00000000001011111000010000101011;
				12'h969: data <= 32'b00000000001011111011001111000111;
				12'h96A: data <= 32'b00000000001011111110001110010011;
				12'h96B: data <= 32'b00000000001100000001001110001110;
				12'h96C: data <= 32'b00000000001100000100001110111010;
				12'h96D: data <= 32'b00000000001100000111010000010110;
				12'h96E: data <= 32'b00000000001100001010010010100010;
				12'h96F: data <= 32'b00000000001100001101010101011111;
				12'h970: data <= 32'b00000000001100010000011001001101;
				12'h971: data <= 32'b00000000001100010011011101101100;
				12'h972: data <= 32'b00000000001100010110100010111100;
				12'h973: data <= 32'b00000000001100011001101000111101;
				12'h974: data <= 32'b00000000001100011100101111110000;
				12'h975: data <= 32'b00000000001100011111110111010101;
				12'h976: data <= 32'b00000000001100100010111111101100;
				12'h977: data <= 32'b00000000001100100110001000110101;
				12'h978: data <= 32'b00000000001100101001010010110000;
				12'h979: data <= 32'b00000000001100101100011101011110;
				12'h97A: data <= 32'b00000000001100101111101000111111;
				12'h97B: data <= 32'b00000000001100110010110101010011;
				12'h97C: data <= 32'b00000000001100110110000010011010;
				12'h97D: data <= 32'b00000000001100111001010000010100;
				12'h97E: data <= 32'b00000000001100111100011111000010;
				12'h97F: data <= 32'b00000000001100111111101110100100;
				12'h980: data <= 32'b00000000001101000010111110111010;
				12'h981: data <= 32'b00000000001101000110010000000011;
				12'h982: data <= 32'b00000000001101001001100010000010;
				12'h983: data <= 32'b00000000001101001100110100110101;
				12'h984: data <= 32'b00000000001101010000001000011100;
				12'h985: data <= 32'b00000000001101010011011100111001;
				12'h986: data <= 32'b00000000001101010110110010001011;
				12'h987: data <= 32'b00000000001101011010001000010010;
				12'h988: data <= 32'b00000000001101011101011111001111;
				12'h989: data <= 32'b00000000001101100000110111000010;
				12'h98A: data <= 32'b00000000001101100100001111101010;
				12'h98B: data <= 32'b00000000001101100111101001001010;
				12'h98C: data <= 32'b00000000001101101011000011011111;
				12'h98D: data <= 32'b00000000001101101110011110101011;
				12'h98E: data <= 32'b00000000001101110001111010101111;
				12'h98F: data <= 32'b00000000001101110101010111101001;
				12'h990: data <= 32'b00000000001101111000110101011010;
				12'h991: data <= 32'b00000000001101111100010100000100;
				12'h992: data <= 32'b00000000001101111111110011100101;
				12'h993: data <= 32'b00000000001110000011010011111101;
				12'h994: data <= 32'b00000000001110000110110101001111;
				12'h995: data <= 32'b00000000001110001010010111011000;
				12'h996: data <= 32'b00000000001110001101111010011010;
				12'h997: data <= 32'b00000000001110010001011110010101;
				12'h998: data <= 32'b00000000001110010101000011001010;
				12'h999: data <= 32'b00000000001110011000101000110111;
				12'h99A: data <= 32'b00000000001110011100001111011110;
				12'h99B: data <= 32'b00000000001110011111110110111111;
				12'h99C: data <= 32'b00000000001110100011011111011010;
				12'h99D: data <= 32'b00000000001110100111001000101111;
				12'h99E: data <= 32'b00000000001110101010110010111110;
				12'h99F: data <= 32'b00000000001110101110011110001000;
				12'h9A0: data <= 32'b00000000001110110010001010001101;
				12'h9A1: data <= 32'b00000000001110110101110111001101;
				12'h9A2: data <= 32'b00000000001110111001100101001001;
				12'h9A3: data <= 32'b00000000001110111101010100000000;
				12'h9A4: data <= 32'b00000000001111000001000011110011;
				12'h9A5: data <= 32'b00000000001111000100110100100010;
				12'h9A6: data <= 32'b00000000001111001000100110001101;
				12'h9A7: data <= 32'b00000000001111001100011000110101;
				12'h9A8: data <= 32'b00000000001111010000001100011010;
				12'h9A9: data <= 32'b00000000001111010100000000111100;
				12'h9AA: data <= 32'b00000000001111010111110110011010;
				12'h9AB: data <= 32'b00000000001111011011101100110111;
				12'h9AC: data <= 32'b00000000001111011111100100010001;
				12'h9AD: data <= 32'b00000000001111100011011100101001;
				12'h9AE: data <= 32'b00000000001111100111010101111111;
				12'h9AF: data <= 32'b00000000001111101011010000010100;
				12'h9B0: data <= 32'b00000000001111101111001011101000;
				12'h9B1: data <= 32'b00000000001111110011000111111010;
				12'h9B2: data <= 32'b00000000001111110111000101001100;
				12'h9B3: data <= 32'b00000000001111111011000011011101;
				12'h9B4: data <= 32'b00000000001111111111000010101101;
				12'h9B5: data <= 32'b00000000010000000011000010111110;
				12'h9B6: data <= 32'b00000000010000000111000100001111;
				12'h9B7: data <= 32'b00000000010000001011000110100000;
				12'h9B8: data <= 32'b00000000010000001111001001110010;
				12'h9B9: data <= 32'b00000000010000010011001110000101;
				12'h9BA: data <= 32'b00000000010000010111010011011001;
				12'h9BB: data <= 32'b00000000010000011011011001101111;
				12'h9BC: data <= 32'b00000000010000011111100001000110;
				12'h9BD: data <= 32'b00000000010000100011101001100000;
				12'h9BE: data <= 32'b00000000010000100111110010111011;
				12'h9BF: data <= 32'b00000000010000101011111101011001;
				12'h9C0: data <= 32'b00000000010000110000001000111010;
				12'h9C1: data <= 32'b00000000010000110100010101011110;
				12'h9C2: data <= 32'b00000000010000111000100011000101;
				12'h9C3: data <= 32'b00000000010000111100110001101111;
				12'h9C4: data <= 32'b00000000010001000001000001011110;
				12'h9C5: data <= 32'b00000000010001000101010010010000;
				12'h9C6: data <= 32'b00000000010001001001100100000111;
				12'h9C7: data <= 32'b00000000010001001101110111000010;
				12'h9C8: data <= 32'b00000000010001010010001011000011;
				12'h9C9: data <= 32'b00000000010001010110100000001000;
				12'h9CA: data <= 32'b00000000010001011010110110010011;
				12'h9CB: data <= 32'b00000000010001011111001101100011;
				12'h9CC: data <= 32'b00000000010001100011100101111010;
				12'h9CD: data <= 32'b00000000010001100111111111010110;
				12'h9CE: data <= 32'b00000000010001101100011001111001;
				12'h9CF: data <= 32'b00000000010001110000110101100011;
				12'h9D0: data <= 32'b00000000010001110101010010010100;
				12'h9D1: data <= 32'b00000000010001111001110000001101;
				12'h9D2: data <= 32'b00000000010001111110001111001101;
				12'h9D3: data <= 32'b00000000010010000010101111010100;
				12'h9D4: data <= 32'b00000000010010000111010000100100;
				12'h9D5: data <= 32'b00000000010010001011110010111101;
				12'h9D6: data <= 32'b00000000010010010000010110011110;
				12'h9D7: data <= 32'b00000000010010010100111011001000;
				12'h9D8: data <= 32'b00000000010010011001100000111100;
				12'h9D9: data <= 32'b00000000010010011110000111111001;
				12'h9DA: data <= 32'b00000000010010100010110000000000;
				12'h9DB: data <= 32'b00000000010010100111011001010001;
				12'h9DC: data <= 32'b00000000010010101100000011101100;
				12'h9DD: data <= 32'b00000000010010110000101111010011;
				12'h9DE: data <= 32'b00000000010010110101011100000100;
				12'h9DF: data <= 32'b00000000010010111010001010000001;
				12'h9E0: data <= 32'b00000000010010111110111001001001;
				12'h9E1: data <= 32'b00000000010011000011101001011101;
				12'h9E2: data <= 32'b00000000010011001000011010111110;
				12'h9E3: data <= 32'b00000000010011001101001101101011;
				12'h9E4: data <= 32'b00000000010011010010000001100101;
				12'h9E5: data <= 32'b00000000010011010110110110101100;
				12'h9E6: data <= 32'b00000000010011011011101101000000;
				12'h9E7: data <= 32'b00000000010011100000100100100011;
				12'h9E8: data <= 32'b00000000010011100101011101010011;
				12'h9E9: data <= 32'b00000000010011101010010111010001;
				12'h9EA: data <= 32'b00000000010011101111010010011111;
				12'h9EB: data <= 32'b00000000010011110100001110111011;
				12'h9EC: data <= 32'b00000000010011111001001100100110;
				12'h9ED: data <= 32'b00000000010011111110001011100001;
				12'h9EE: data <= 32'b00000000010100000011001011101100;
				12'h9EF: data <= 32'b00000000010100001000001101000111;
				12'h9F0: data <= 32'b00000000010100001101001111110011;
				12'h9F1: data <= 32'b00000000010100010010010011101111;
				12'h9F2: data <= 32'b00000000010100010111011000111101;
				12'h9F3: data <= 32'b00000000010100011100011111011100;
				12'h9F4: data <= 32'b00000000010100100001100111001100;
				12'h9F5: data <= 32'b00000000010100100110110000001111;
				12'h9F6: data <= 32'b00000000010100101011111010100101;
				12'h9F7: data <= 32'b00000000010100110001000110001101;
				12'h9F8: data <= 32'b00000000010100110110010011001000;
				12'h9F9: data <= 32'b00000000010100111011100001010110;
				12'h9FA: data <= 32'b00000000010101000000110000111001;
				12'h9FB: data <= 32'b00000000010101000110000001101111;
				12'h9FC: data <= 32'b00000000010101001011010011111010;
				12'h9FD: data <= 32'b00000000010101010000100111011001;
				12'h9FE: data <= 32'b00000000010101010101111100001101;
				12'h9FF: data <= 32'b00000000010101011011010010010111;
				12'hA00: data <= 32'b00000000010101100000101001110111;
				12'hA01: data <= 32'b00000000010101100110000010101100;
				12'hA02: data <= 32'b00000000010101101011011100111000;
				12'hA03: data <= 32'b00000000010101110000111000011011;
				12'hA04: data <= 32'b00000000010101110110010101010101;
				12'hA05: data <= 32'b00000000010101111011110011100110;
				12'hA06: data <= 32'b00000000010110000001010011001110;
				12'hA07: data <= 32'b00000000010110000110110100001111;
				12'hA08: data <= 32'b00000000010110001100010110101001;
				12'hA09: data <= 32'b00000000010110010001111010011011;
				12'hA0A: data <= 32'b00000000010110010111011111100110;
				12'hA0B: data <= 32'b00000000010110011101000110001011;
				12'hA0C: data <= 32'b00000000010110100010101110001001;
				12'hA0D: data <= 32'b00000000010110101000010111100010;
				12'hA0E: data <= 32'b00000000010110101110000010010101;
				12'hA0F: data <= 32'b00000000010110110011101110100011;
				12'hA10: data <= 32'b00000000010110111001011100001101;
				12'hA11: data <= 32'b00000000010110111111001011010001;
				12'hA12: data <= 32'b00000000010111000100111011110010;
				12'hA13: data <= 32'b00000000010111001010101101101111;
				12'hA14: data <= 32'b00000000010111010000100001001001;
				12'hA15: data <= 32'b00000000010111010110010110000000;
				12'hA16: data <= 32'b00000000010111011100001100010100;
				12'hA17: data <= 32'b00000000010111100010000100000110;
				12'hA18: data <= 32'b00000000010111100111111101010111;
				12'hA19: data <= 32'b00000000010111101101111000000101;
				12'hA1A: data <= 32'b00000000010111110011110100010011;
				12'hA1B: data <= 32'b00000000010111111001110001111111;
				12'hA1C: data <= 32'b00000000010111111111110001001100;
				12'hA1D: data <= 32'b00000000011000000101110001111000;
				12'hA1E: data <= 32'b00000000011000001011110100000101;
				12'hA1F: data <= 32'b00000000011000010001110111110010;
				12'hA20: data <= 32'b00000000011000010111111101000001;
				12'hA21: data <= 32'b00000000011000011110000011110001;
				12'hA22: data <= 32'b00000000011000100100001100000011;
				12'hA23: data <= 32'b00000000011000101010010101110111;
				12'hA24: data <= 32'b00000000011000110000100001001110;
				12'hA25: data <= 32'b00000000011000110110101110001000;
				12'hA26: data <= 32'b00000000011000111100111100100101;
				12'hA27: data <= 32'b00000000011001000011001100100110;
				12'hA28: data <= 32'b00000000011001001001011110001100;
				12'hA29: data <= 32'b00000000011001001111110001010110;
				12'hA2A: data <= 32'b00000000011001010110000110000100;
				12'hA2B: data <= 32'b00000000011001011100011100011001;
				12'hA2C: data <= 32'b00000000011001100010110100010011;
				12'hA2D: data <= 32'b00000000011001101001001101110011;
				12'hA2E: data <= 32'b00000000011001101111101000111010;
				12'hA2F: data <= 32'b00000000011001110110000101101000;
				12'hA30: data <= 32'b00000000011001111100100011111101;
				12'hA31: data <= 32'b00000000011010000011000011111010;
				12'hA32: data <= 32'b00000000011010001001100101011111;
				12'hA33: data <= 32'b00000000011010010000001000101101;
				12'hA34: data <= 32'b00000000011010010110101101100011;
				12'hA35: data <= 32'b00000000011010011101010100000100;
				12'hA36: data <= 32'b00000000011010100011111100001110;
				12'hA37: data <= 32'b00000000011010101010100110000010;
				12'hA38: data <= 32'b00000000011010110001010001100001;
				12'hA39: data <= 32'b00000000011010110111111110101011;
				12'hA3A: data <= 32'b00000000011010111110101101100000;
				12'hA3B: data <= 32'b00000000011011000101011110000010;
				12'hA3C: data <= 32'b00000000011011001100010000001111;
				12'hA3D: data <= 32'b00000000011011010011000100001010;
				12'hA3E: data <= 32'b00000000011011011001111001110010;
				12'hA3F: data <= 32'b00000000011011100000110001000111;
				12'hA40: data <= 32'b00000000011011100111101010001010;
				12'hA41: data <= 32'b00000000011011101110100100111100;
				12'hA42: data <= 32'b00000000011011110101100001011101;
				12'hA43: data <= 32'b00000000011011111100011111101101;
				12'hA44: data <= 32'b00000000011100000011011111101101;
				12'hA45: data <= 32'b00000000011100001010100001011101;
				12'hA46: data <= 32'b00000000011100010001100100111110;
				12'hA47: data <= 32'b00000000011100011000101010010000;
				12'hA48: data <= 32'b00000000011100011111110001010011;
				12'hA49: data <= 32'b00000000011100100110111010001000;
				12'hA4A: data <= 32'b00000000011100101110000100110000;
				12'hA4B: data <= 32'b00000000011100110101010001001011;
				12'hA4C: data <= 32'b00000000011100111100011111011001;
				12'hA4D: data <= 32'b00000000011101000011101111011011;
				12'hA4E: data <= 32'b00000000011101001011000001010001;
				12'hA4F: data <= 32'b00000000011101010010010100111100;
				12'hA50: data <= 32'b00000000011101011001101010011011;
				12'hA51: data <= 32'b00000000011101100001000001110001;
				12'hA52: data <= 32'b00000000011101101000011010111100;
				12'hA53: data <= 32'b00000000011101101111110101111111;
				12'hA54: data <= 32'b00000000011101110111010010111000;
				12'hA55: data <= 32'b00000000011101111110110001101000;
				12'hA56: data <= 32'b00000000011110000110010010010001;
				12'hA57: data <= 32'b00000000011110001101110100110001;
				12'hA58: data <= 32'b00000000011110010101011001001011;
				12'hA59: data <= 32'b00000000011110011100111111011110;
				12'hA5A: data <= 32'b00000000011110100100100111101011;
				12'hA5B: data <= 32'b00000000011110101100010001110010;
				12'hA5C: data <= 32'b00000000011110110011111101110100;
				12'hA5D: data <= 32'b00000000011110111011101011110001;
				12'hA5E: data <= 32'b00000000011111000011011011101010;
				12'hA5F: data <= 32'b00000000011111001011001101011111;
				12'hA60: data <= 32'b00000000011111010011000001010001;
				12'hA61: data <= 32'b00000000011111011010110111000000;
				12'hA62: data <= 32'b00000000011111100010101110101101;
				12'hA63: data <= 32'b00000000011111101010101000011000;
				12'hA64: data <= 32'b00000000011111110010100100000001;
				12'hA65: data <= 32'b00000000011111111010100001101010;
				12'hA66: data <= 32'b00000000100000000010100001010010;
				12'hA67: data <= 32'b00000000100000001010100010111011;
				12'hA68: data <= 32'b00000000100000010010100110100100;
				12'hA69: data <= 32'b00000000100000011010101100001110;
				12'hA6A: data <= 32'b00000000100000100010110011111010;
				12'hA6B: data <= 32'b00000000100000101010111101101000;
				12'hA6C: data <= 32'b00000000100000110011001001011001;
				12'hA6D: data <= 32'b00000000100000111011010111001101;
				12'hA6E: data <= 32'b00000000100001000011100111000101;
				12'hA6F: data <= 32'b00000000100001001011111001000001;
				12'hA70: data <= 32'b00000000100001010100001101000001;
				12'hA71: data <= 32'b00000000100001011100100011000111;
				12'hA72: data <= 32'b00000000100001100100111011010011;
				12'hA73: data <= 32'b00000000100001101101010101100101;
				12'hA74: data <= 32'b00000000100001110101110001111110;
				12'hA75: data <= 32'b00000000100001111110010000011110;
				12'hA76: data <= 32'b00000000100010000110110001000111;
				12'hA77: data <= 32'b00000000100010001111010011110111;
				12'hA78: data <= 32'b00000000100010010111111000110001;
				12'hA79: data <= 32'b00000000100010100000011111110100;
				12'hA7A: data <= 32'b00000000100010101001001001000001;
				12'hA7B: data <= 32'b00000000100010110001110100011000;
				12'hA7C: data <= 32'b00000000100010111010100001111011;
				12'hA7D: data <= 32'b00000000100011000011010001101010;
				12'hA7E: data <= 32'b00000000100011001100000011100100;
				12'hA7F: data <= 32'b00000000100011010100110111101100;
				12'hA80: data <= 32'b00000000100011011101101110000000;
				12'hA81: data <= 32'b00000000100011100110100110100011;
				12'hA82: data <= 32'b00000000100011101111100001010100;
				12'hA83: data <= 32'b00000000100011111000011110010100;
				12'hA84: data <= 32'b00000000100100000001011101100011;
				12'hA85: data <= 32'b00000000100100001010011111000011;
				12'hA86: data <= 32'b00000000100100010011100010110011;
				12'hA87: data <= 32'b00000000100100011100101000110100;
				12'hA88: data <= 32'b00000000100100100101110001000111;
				12'hA89: data <= 32'b00000000100100101110111011101101;
				12'hA8A: data <= 32'b00000000100100111000001000100101;
				12'hA8B: data <= 32'b00000000100101000001010111110001;
				12'hA8C: data <= 32'b00000000100101001010101001010001;
				12'hA8D: data <= 32'b00000000100101010011111101000110;
				12'hA8E: data <= 32'b00000000100101011101010011010000;
				12'hA8F: data <= 32'b00000000100101100110101011110000;
				12'hA90: data <= 32'b00000000100101110000000110100110;
				12'hA91: data <= 32'b00000000100101111001100011110100;
				12'hA92: data <= 32'b00000000100110000011000011011000;
				12'hA93: data <= 32'b00000000100110001100100101010101;
				12'hA94: data <= 32'b00000000100110010110001001101011;
				12'hA95: data <= 32'b00000000100110011111110000011010;
				12'hA96: data <= 32'b00000000100110101001011001100100;
				12'hA97: data <= 32'b00000000100110110011000101000111;
				12'hA98: data <= 32'b00000000100110111100110011000110;
				12'hA99: data <= 32'b00000000100111000110100011100001;
				12'hA9A: data <= 32'b00000000100111010000010110011000;
				12'hA9B: data <= 32'b00000000100111011010001011101101;
				12'hA9C: data <= 32'b00000000100111100100000011011110;
				12'hA9D: data <= 32'b00000000100111101101111101101111;
				12'hA9E: data <= 32'b00000000100111110111111010011101;
				12'hA9F: data <= 32'b00000000101000000001111001101100;
				12'hAA0: data <= 32'b00000000101000001011111011011011;
				12'hAA1: data <= 32'b00000000101000010101111111101010;
				12'hAA2: data <= 32'b00000000101000100000000110011011;
				12'hAA3: data <= 32'b00000000101000101010001111101101;
				12'hAA4: data <= 32'b00000000101000110100011011100011;
				12'hAA5: data <= 32'b00000000101000111110101001111011;
				12'hAA6: data <= 32'b00000000101001001000111010111000;
				12'hAA7: data <= 32'b00000000101001010011001110011001;
				12'hAA8: data <= 32'b00000000101001011101100100011111;
				12'hAA9: data <= 32'b00000000101001100111111101001011;
				12'hAAA: data <= 32'b00000000101001110010011000011110;
				12'hAAB: data <= 32'b00000000101001111100110110011000;
				12'hAAC: data <= 32'b00000000101010000111010110111001;
				12'hAAD: data <= 32'b00000000101010010001111010000100;
				12'hAAE: data <= 32'b00000000101010011100011111110111;
				12'hAAF: data <= 32'b00000000101010100111001000010100;
				12'hAB0: data <= 32'b00000000101010110001110011011011;
				12'hAB1: data <= 32'b00000000101010111100100001001110;
				12'hAB2: data <= 32'b00000000101011000111010001101100;
				12'hAB3: data <= 32'b00000000101011010010000100110111;
				12'hAB4: data <= 32'b00000000101011011100111010101111;
				12'hAB5: data <= 32'b00000000101011100111110011010100;
				12'hAB6: data <= 32'b00000000101011110010101110101000;
				12'hAB7: data <= 32'b00000000101011111101101100101100;
				12'hAB8: data <= 32'b00000000101100001000101101011111;
				12'hAB9: data <= 32'b00000000101100010011110001000011;
				12'hABA: data <= 32'b00000000101100011110110111011000;
				12'hABB: data <= 32'b00000000101100101010000000011111;
				12'hABC: data <= 32'b00000000101100110101001100011000;
				12'hABD: data <= 32'b00000000101101000000011011000101;
				12'hABE: data <= 32'b00000000101101001011101100100110;
				12'hABF: data <= 32'b00000000101101010111000000111100;
				12'hAC0: data <= 32'b00000000101101100010011000000111;
				12'hAC1: data <= 32'b00000000101101101101110010001000;
				12'hAC2: data <= 32'b00000000101101111001001111000000;
				12'hAC3: data <= 32'b00000000101110000100101110110000;
				12'hAC4: data <= 32'b00000000101110010000010001011000;
				12'hAC5: data <= 32'b00000000101110011011110110111001;
				12'hAC6: data <= 32'b00000000101110100111011111010011;
				12'hAC7: data <= 32'b00000000101110110011001010101001;
				12'hAC8: data <= 32'b00000000101110111110111000111001;
				12'hAC9: data <= 32'b00000000101111001010101010000101;
				12'hACA: data <= 32'b00000000101111010110011110001110;
				12'hACB: data <= 32'b00000000101111100010010101010101;
				12'hACC: data <= 32'b00000000101111101110001111011001;
				12'hACD: data <= 32'b00000000101111111010001100011101;
				12'hACE: data <= 32'b00000000110000000110001100100000;
				12'hACF: data <= 32'b00000000110000010010001111100011;
				12'hAD0: data <= 32'b00000000110000011110010101101000;
				12'hAD1: data <= 32'b00000000110000101010011110101110;
				12'hAD2: data <= 32'b00000000110000110110101010110111;
				12'hAD3: data <= 32'b00000000110001000010111010000100;
				12'hAD4: data <= 32'b00000000110001001111001100010101;
				12'hAD5: data <= 32'b00000000110001011011100001101010;
				12'hAD6: data <= 32'b00000000110001100111111010000110;
				12'hAD7: data <= 32'b00000000110001110100010101101000;
				12'hAD8: data <= 32'b00000000110010000000110100010001;
				12'hAD9: data <= 32'b00000000110010001101010110000010;
				12'hADA: data <= 32'b00000000110010011001111010111100;
				12'hADB: data <= 32'b00000000110010100110100011000000;
				12'hADC: data <= 32'b00000000110010110011001110001110;
				12'hADD: data <= 32'b00000000110010111111111100100111;
				12'hADE: data <= 32'b00000000110011001100101110001100;
				12'hADF: data <= 32'b00000000110011011001100010111110;
				12'hAE0: data <= 32'b00000000110011100110011010111110;
				12'hAE1: data <= 32'b00000000110011110011010110001100;
				12'hAE2: data <= 32'b00000000110100000000010100101001;
				12'hAE3: data <= 32'b00000000110100001101010110010111;
				12'hAE4: data <= 32'b00000000110100011010011011010101;
				12'hAE5: data <= 32'b00000000110100100111100011100101;
				12'hAE6: data <= 32'b00000000110100110100101111000111;
				12'hAE7: data <= 32'b00000000110101000001111101111101;
				12'hAE8: data <= 32'b00000000110101001111010000000110;
				12'hAE9: data <= 32'b00000000110101011100100101100101;
				12'hAEA: data <= 32'b00000000110101101001111110011001;
				12'hAEB: data <= 32'b00000000110101110111011010100100;
				12'hAEC: data <= 32'b00000000110110000100111010000111;
				12'hAED: data <= 32'b00000000110110010010011101000010;
				12'hAEE: data <= 32'b00000000110110100000000011010110;
				12'hAEF: data <= 32'b00000000110110101101101101000100;
				12'hAF0: data <= 32'b00000000110110111011011010001101;
				12'hAF1: data <= 32'b00000000110111001001001010110001;
				12'hAF2: data <= 32'b00000000110111010110111110110010;
				12'hAF3: data <= 32'b00000000110111100100110110010001;
				12'hAF4: data <= 32'b00000000110111110010110001001110;
				12'hAF5: data <= 32'b00000000111000000000101111101010;
				12'hAF6: data <= 32'b00000000111000001110110001100110;
				12'hAF7: data <= 32'b00000000111000011100110111000011;
				12'hAF8: data <= 32'b00000000111000101011000000000010;
				12'hAF9: data <= 32'b00000000111000111001001100100011;
				12'hAFA: data <= 32'b00000000111001000111011100101000;
				12'hAFB: data <= 32'b00000000111001010101110000010010;
				12'hAFC: data <= 32'b00000000111001100100000111100001;
				12'hAFD: data <= 32'b00000000111001110010100010010110;
				12'hAFE: data <= 32'b00000000111010000001000000110010;
				12'hAFF: data <= 32'b00000000111010001111100010110110;
				12'hB00: data <= 32'b00000000111010011110001000100100;
				12'hB01: data <= 32'b00000000111010101100110001111011;
				12'hB02: data <= 32'b00000000111010111011011110111101;
				12'hB03: data <= 32'b00000000111011001010001111101011;
				12'hB04: data <= 32'b00000000111011011001000100000101;
				12'hB05: data <= 32'b00000000111011100111111100001101;
				12'hB06: data <= 32'b00000000111011110110111000000100;
				12'hB07: data <= 32'b00000000111100000101110111101010;
				12'hB08: data <= 32'b00000000111100010100111011000000;
				12'hB09: data <= 32'b00000000111100100100000010000111;
				12'hB0A: data <= 32'b00000000111100110011001101000001;
				12'hB0B: data <= 32'b00000000111101000010011011101110;
				12'hB0C: data <= 32'b00000000111101010001101110001111;
				12'hB0D: data <= 32'b00000000111101100001000100100110;
				12'hB0E: data <= 32'b00000000111101110000011110110010;
				12'hB0F: data <= 32'b00000000111101111111111100110101;
				12'hB10: data <= 32'b00000000111110001111011110110001;
				12'hB11: data <= 32'b00000000111110011111000100100101;
				12'hB12: data <= 32'b00000000111110101110101110010011;
				12'hB13: data <= 32'b00000000111110111110011011111100;
				12'hB14: data <= 32'b00000000111111001110001101100010;
				12'hB15: data <= 32'b00000000111111011110000011000100;
				12'hB16: data <= 32'b00000000111111101101111100100011;
				12'hB17: data <= 32'b00000000111111111101111010000010;
				12'hB18: data <= 32'b00000001000000001101111011100001;
				12'hB19: data <= 32'b00000001000000011110000001000000;
				12'hB1A: data <= 32'b00000001000000101110001010100010;
				12'hB1B: data <= 32'b00000001000000111110011000000110;
				12'hB1C: data <= 32'b00000001000001001110101001101110;
				12'hB1D: data <= 32'b00000001000001011110111111011011;
				12'hB1E: data <= 32'b00000001000001101111011001001110;
				12'hB1F: data <= 32'b00000001000001111111110111001000;
				12'hB20: data <= 32'b00000001000010010000011001001010;
				12'hB21: data <= 32'b00000001000010100000111111010101;
				12'hB22: data <= 32'b00000001000010110001101001101010;
				12'hB23: data <= 32'b00000001000011000010011000001010;
				12'hB24: data <= 32'b00000001000011010011001010110110;
				12'hB25: data <= 32'b00000001000011100100000001110000;
				12'hB26: data <= 32'b00000001000011110100111100111000;
				12'hB27: data <= 32'b00000001000100000101111100001111;
				12'hB28: data <= 32'b00000001000100010110111111110110;
				12'hB29: data <= 32'b00000001000100101000000111101111;
				12'hB2A: data <= 32'b00000001000100111001010011111010;
				12'hB2B: data <= 32'b00000001000101001010100100011001;
				12'hB2C: data <= 32'b00000001000101011011111001001101;
				12'hB2D: data <= 32'b00000001000101101101010010010110;
				12'hB2E: data <= 32'b00000001000101111110101111110110;
				12'hB2F: data <= 32'b00000001000110010000010001101111;
				12'hB30: data <= 32'b00000001000110100001111000000000;
				12'hB31: data <= 32'b00000001000110110011100010101011;
				12'hB32: data <= 32'b00000001000111000101010001110001;
				12'hB33: data <= 32'b00000001000111010111000101010100;
				12'hB34: data <= 32'b00000001000111101000111101010100;
				12'hB35: data <= 32'b00000001000111111010111001110011;
				12'hB36: data <= 32'b00000001001000001100111010110010;
				12'hB37: data <= 32'b00000001001000011111000000010001;
				12'hB38: data <= 32'b00000001001000110001001010010010;
				12'hB39: data <= 32'b00000001001001000011011000110111;
				12'hB3A: data <= 32'b00000001001001010101101011111111;
				12'hB3B: data <= 32'b00000001001001101000000011101101;
				12'hB3C: data <= 32'b00000001001001111010100000000001;
				12'hB3D: data <= 32'b00000001001010001101000000111101;
				12'hB3E: data <= 32'b00000001001010011111100110100010;
				12'hB3F: data <= 32'b00000001001010110010010000110001;
				12'hB40: data <= 32'b00000001001011000100111111101011;
				12'hB41: data <= 32'b00000001001011010111110011010001;
				12'hB42: data <= 32'b00000001001011101010101011100101;
				12'hB43: data <= 32'b00000001001011111101101000100111;
				12'hB44: data <= 32'b00000001001100010000101010011010;
				12'hB45: data <= 32'b00000001001100100011110000111101;
				12'hB46: data <= 32'b00000001001100110110111100010011;
				12'hB47: data <= 32'b00000001001101001010001100011100;
				12'hB48: data <= 32'b00000001001101011101100001011001;
				12'hB49: data <= 32'b00000001001101110000111011001101;
				12'hB4A: data <= 32'b00000001001110000100011001110111;
				12'hB4B: data <= 32'b00000001001110010111111101011010;
				12'hB4C: data <= 32'b00000001001110101011100101110110;
				12'hB4D: data <= 32'b00000001001110111111010011001101;
				12'hB4E: data <= 32'b00000001001111010011000101100000;
				12'hB4F: data <= 32'b00000001001111100110111100110001;
				12'hB50: data <= 32'b00000001001111111010111000111111;
				12'hB51: data <= 32'b00000001010000001110111010001101;
				12'hB52: data <= 32'b00000001010000100011000000011101;
				12'hB53: data <= 32'b00000001010000110111001011101110;
				12'hB54: data <= 32'b00000001010001001011011100000011;
				12'hB55: data <= 32'b00000001010001011111110001011101;
				12'hB56: data <= 32'b00000001010001110100001011111100;
				12'hB57: data <= 32'b00000001010010001000101011100011;
				12'hB58: data <= 32'b00000001010010011101010000010010;
				12'hB59: data <= 32'b00000001010010110001111010001100;
				12'hB5A: data <= 32'b00000001010011000110101001010000;
				12'hB5B: data <= 32'b00000001010011011011011101100001;
				12'hB5C: data <= 32'b00000001010011110000010110111111;
				12'hB5D: data <= 32'b00000001010100000101010101101101;
				12'hB5E: data <= 32'b00000001010100011010011001101010;
				12'hB5F: data <= 32'b00000001010100101111100010111010;
				12'hB60: data <= 32'b00000001010101000100110001011100;
				12'hB61: data <= 32'b00000001010101011010000101010011;
				12'hB62: data <= 32'b00000001010101101111011110011111;
				12'hB63: data <= 32'b00000001010110000100111101000011;
				12'hB64: data <= 32'b00000001010110011010100000111110;
				12'hB65: data <= 32'b00000001010110110000001010010100;
				12'hB66: data <= 32'b00000001010111000101111001000100;
				12'hB67: data <= 32'b00000001010111011011101101010001;
				12'hB68: data <= 32'b00000001010111110001100110111011;
				12'hB69: data <= 32'b00000001011000000111100110000100;
				12'hB6A: data <= 32'b00000001011000011101101010101110;
				12'hB6B: data <= 32'b00000001011000110011110100111010;
				12'hB6C: data <= 32'b00000001011001001010000100101001;
				12'hB6D: data <= 32'b00000001011001100000011001111101;
				12'hB6E: data <= 32'b00000001011001110110110100110111;
				12'hB6F: data <= 32'b00000001011010001101010101011000;
				12'hB70: data <= 32'b00000001011010100011111011100010;
				12'hB71: data <= 32'b00000001011010111010100111010110;
				12'hB72: data <= 32'b00000001011011010001011000110110;
				12'hB73: data <= 32'b00000001011011101000010000000011;
				12'hB74: data <= 32'b00000001011011111111001100111111;
				12'hB75: data <= 32'b00000001011100010110001111101010;
				12'hB76: data <= 32'b00000001011100101101011000000111;
				12'hB77: data <= 32'b00000001011101000100100110010111;
				12'hB78: data <= 32'b00000001011101011011111010011011;
				12'hB79: data <= 32'b00000001011101110011010100010100;
				12'hB7A: data <= 32'b00000001011110001010110100000101;
				12'hB7B: data <= 32'b00000001011110100010011001101111;
				12'hB7C: data <= 32'b00000001011110111010000101010011;
				12'hB7D: data <= 32'b00000001011111010001110110110010;
				12'hB7E: data <= 32'b00000001011111101001101110001111;
				12'hB7F: data <= 32'b00000001100000000001101011101010;
				12'hB80: data <= 32'b00000001100000011001101111000101;
				12'hB81: data <= 32'b00000001100000110001111000100010;
				12'hB82: data <= 32'b00000001100001001010001000000010;
				12'hB83: data <= 32'b00000001100001100010011101100110;
				12'hB84: data <= 32'b00000001100001111010111001010001;
				12'hB85: data <= 32'b00000001100010010011011011000011;
				12'hB86: data <= 32'b00000001100010101100000010111111;
				12'hB87: data <= 32'b00000001100011000100110001000101;
				12'hB88: data <= 32'b00000001100011011101100101011000;
				12'hB89: data <= 32'b00000001100011110110011111111001;
				12'hB8A: data <= 32'b00000001100100001111100000101001;
				12'hB8B: data <= 32'b00000001100100101000100111101001;
				12'hB8C: data <= 32'b00000001100101000001110100111101;
				12'hB8D: data <= 32'b00000001100101011011001000100100;
				12'hB8E: data <= 32'b00000001100101110100100010100010;
				12'hB8F: data <= 32'b00000001100110001110000010110110;
				12'hB90: data <= 32'b00000001100110100111101001100100;
				12'hB91: data <= 32'b00000001100111000001010110101100;
				12'hB92: data <= 32'b00000001100111011011001010010000;
				12'hB93: data <= 32'b00000001100111110101000100010001;
				12'hB94: data <= 32'b00000001101000001111000100110010;
				12'hB95: data <= 32'b00000001101000101001001011110100;
				12'hB96: data <= 32'b00000001101001000011011001011001;
				12'hB97: data <= 32'b00000001101001011101101101100001;
				12'hB98: data <= 32'b00000001101001111000001000010000;
				12'hB99: data <= 32'b00000001101010010010101001100110;
				12'hB9A: data <= 32'b00000001101010101101010001100101;
				12'hB9B: data <= 32'b00000001101011001000000000001111;
				12'hB9C: data <= 32'b00000001101011100010110101100110;
				12'hB9D: data <= 32'b00000001101011111101110001101011;
				12'hB9E: data <= 32'b00000001101100011000110100011111;
				12'hB9F: data <= 32'b00000001101100110011111110000110;
				12'hBA0: data <= 32'b00000001101101001111001110011111;
				12'hBA1: data <= 32'b00000001101101101010100101101101;
				12'hBA2: data <= 32'b00000001101110000110000011110010;
				12'hBA3: data <= 32'b00000001101110100001101000110000;
				12'hBA4: data <= 32'b00000001101110111101010100100111;
				12'hBA5: data <= 32'b00000001101111011001000111011011;
				12'hBA6: data <= 32'b00000001101111110101000001001100;
				12'hBA7: data <= 32'b00000001110000010001000001111100;
				12'hBA8: data <= 32'b00000001110000101101001001101101;
				12'hBA9: data <= 32'b00000001110001001001011000100001;
				12'hBAA: data <= 32'b00000001110001100101101110011010;
				12'hBAB: data <= 32'b00000001110010000010001011011001;
				12'hBAC: data <= 32'b00000001110010011110101111100000;
				12'hBAD: data <= 32'b00000001110010111011011010110010;
				12'hBAE: data <= 32'b00000001110011011000001101001110;
				12'hBAF: data <= 32'b00000001110011110101000110111001;
				12'hBB0: data <= 32'b00000001110100010010000111110010;
				12'hBB1: data <= 32'b00000001110100101111001111111101;
				12'hBB2: data <= 32'b00000001110101001100011111011011;
				12'hBB3: data <= 32'b00000001110101101001110110001110;
				12'hBB4: data <= 32'b00000001110110000111010100010111;
				12'hBB5: data <= 32'b00000001110110100100111001111000;
				12'hBB6: data <= 32'b00000001110111000010100110110100;
				12'hBB7: data <= 32'b00000001110111100000011011001100;
				12'hBB8: data <= 32'b00000001110111111110010111000011;
				12'hBB9: data <= 32'b00000001111000011100011010011001;
				12'hBBA: data <= 32'b00000001111000111010100101010000;
				12'hBBB: data <= 32'b00000001111001011000110111101100;
				12'hBBC: data <= 32'b00000001111001110111010001101101;
				12'hBBD: data <= 32'b00000001111010010101110011010101;
				12'hBBE: data <= 32'b00000001111010110100011100100111;
				12'hBBF: data <= 32'b00000001111011010011001101100100;
				12'hBC0: data <= 32'b00000001111011110010000110001111;
				12'hBC1: data <= 32'b00000001111100010001000110101000;
				12'hBC2: data <= 32'b00000001111100110000001110110011;
				12'hBC3: data <= 32'b00000001111101001111011110110000;
				12'hBC4: data <= 32'b00000001111101101110110110100011;
				12'hBC5: data <= 32'b00000001111110001110010110001100;
				12'hBC6: data <= 32'b00000001111110101101111101101110;
				12'hBC7: data <= 32'b00000001111111001101101101001100;
				12'hBC8: data <= 32'b00000001111111101101100100100110;
				12'hBC9: data <= 32'b00000010000000001101100011111111;
				12'hBCA: data <= 32'b00000010000000101101101011011000;
				12'hBCB: data <= 32'b00000010000001001101111010110101;
				12'hBCC: data <= 32'b00000010000001101110010010010110;
				12'hBCD: data <= 32'b00000010000010001110110001111111;
				12'hBCE: data <= 32'b00000010000010101111011001110000;
				12'hBCF: data <= 32'b00000010000011010000001001101100;
				12'hBD0: data <= 32'b00000010000011110001000001110110;
				12'hBD1: data <= 32'b00000010000100010010000010001110;
				12'hBD2: data <= 32'b00000010000100110011001010110111;
				12'hBD3: data <= 32'b00000010000101010100011011110100;
				12'hBD4: data <= 32'b00000010000101110101110101000110;
				12'hBD5: data <= 32'b00000010000110010111010110101111;
				12'hBD6: data <= 32'b00000010000110111001000000110010;
				12'hBD7: data <= 32'b00000010000111011010110011010000;
				12'hBD8: data <= 32'b00000010000111111100101110001100;
				12'hBD9: data <= 32'b00000010001000011110110001101000;
				12'hBDA: data <= 32'b00000010001001000000111101100110;
				12'hBDB: data <= 32'b00000010001001100011010010001000;
				12'hBDC: data <= 32'b00000010001010000101101111010000;
				12'hBDD: data <= 32'b00000010001010101000010101000000;
				12'hBDE: data <= 32'b00000010001011001011000011011011;
				12'hBDF: data <= 32'b00000010001011101101111010100010;
				12'hBE0: data <= 32'b00000010001100010000111010011001;
				12'hBE1: data <= 32'b00000010001100110100000011000000;
				12'hBE2: data <= 32'b00000010001101010111010100011011;
				12'hBE3: data <= 32'b00000010001101111010101110101011;
				12'hBE4: data <= 32'b00000010001110011110010001110011;
				12'hBE5: data <= 32'b00000010001111000001111101110101;
				12'hBE6: data <= 32'b00000010001111100101110010110011;
				12'hBE7: data <= 32'b00000010010000001001110000101111;
				12'hBE8: data <= 32'b00000010010000101101110111101100;
				12'hBE9: data <= 32'b00000010010001010010000111101100;
				12'hBEA: data <= 32'b00000010010001110110100000110001;
				12'hBEB: data <= 32'b00000010010010011011000010111101;
				12'hBEC: data <= 32'b00000010010010111111101110010011;
				12'hBED: data <= 32'b00000010010011100100100010110101;
				12'hBEE: data <= 32'b00000010010100001001100000100101;
				12'hBEF: data <= 32'b00000010010100101110100111100110;
				12'hBF0: data <= 32'b00000010010101010011110111111010;
				12'hBF1: data <= 32'b00000010010101111001010001100011;
				12'hBF2: data <= 32'b00000010010110011110110100100011;
				12'hBF3: data <= 32'b00000010010111000100100000111110;
				12'hBF4: data <= 32'b00000010010111101010010110110100;
				12'hBF5: data <= 32'b00000010011000010000010110001010;
				12'hBF6: data <= 32'b00000010011000110110011111000000;
				12'hBF7: data <= 32'b00000010011001011100110001011010;
				12'hBF8: data <= 32'b00000010011010000011001101011010;
				12'hBF9: data <= 32'b00000010011010101001110011000010;
				12'hBFA: data <= 32'b00000010011011010000100010010100;
				12'hBFB: data <= 32'b00000010011011110111011011010100;
				12'hBFC: data <= 32'b00000010011100011110011110000011;
				12'hBFD: data <= 32'b00000010011101000101101010100100;
				12'hBFE: data <= 32'b00000010011101101101000000111001;
				12'hBFF: data <= 32'b00000010011110010100100001000101;
				12'hC00: data <= 32'b00000010011110111100001011001010;
				12'hC01: data <= 32'b00000010011111100011111111001011;
				12'hC02: data <= 32'b00000010100000001011111101001011;
				12'hC03: data <= 32'b00000010100000110100000101001011;
				12'hC04: data <= 32'b00000010100001011100010111001110;
				12'hC05: data <= 32'b00000010100010000100110011010111;
				12'hC06: data <= 32'b00000010100010101101011001101000;
				12'hC07: data <= 32'b00000010100011010110001010000101;
				12'hC08: data <= 32'b00000010100011111111000100101110;
				12'hC09: data <= 32'b00000010100100101000001001101000;
				12'hC0A: data <= 32'b00000010100101010001011000110100;
				12'hC0B: data <= 32'b00000010100101111010110010010101;
				12'hC0C: data <= 32'b00000010100110100100010110001110;
				12'hC0D: data <= 32'b00000010100111001110000100100001;
				12'hC0E: data <= 32'b00000010100111110111111101010001;
				12'hC0F: data <= 32'b00000010101000100010000000100001;
				12'hC10: data <= 32'b00000010101001001100001110010010;
				12'hC11: data <= 32'b00000010101001110110100110101001;
				12'hC12: data <= 32'b00000010101010100001001001100111;
				12'hC13: data <= 32'b00000010101011001011110111001110;
				12'hC14: data <= 32'b00000010101011110110101111100011;
				12'hC15: data <= 32'b00000010101100100001110010100111;
				12'hC16: data <= 32'b00000010101101001101000000011101;
				12'hC17: data <= 32'b00000010101101111000011001001000;
				12'hC18: data <= 32'b00000010101110100011111100101011;
				12'hC19: data <= 32'b00000010101111001111101011000111;
				12'hC1A: data <= 32'b00000010101111111011100100100001;
				12'hC1B: data <= 32'b00000010110000100111101000111011;
				12'hC1C: data <= 32'b00000010110001010011111000010111;
				12'hC1D: data <= 32'b00000010110010000000010010111000;
				12'hC1E: data <= 32'b00000010110010101100111000100001;
				12'hC1F: data <= 32'b00000010110011011001101001010101;
				12'hC20: data <= 32'b00000010110100000110100101010111;
				12'hC21: data <= 32'b00000010110100110011101100101001;
				12'hC22: data <= 32'b00000010110101100000111111001110;
				12'hC23: data <= 32'b00000010110110001110011101001001;
				12'hC24: data <= 32'b00000010110110111100000110011101;
				12'hC25: data <= 32'b00000010110111101001111011001101;
				12'hC26: data <= 32'b00000010111000010111111011011100;
				12'hC27: data <= 32'b00000010111001000110000111001100;
				12'hC28: data <= 32'b00000010111001110100011110100000;
				12'hC29: data <= 32'b00000010111010100011000001011100;
				12'hC2A: data <= 32'b00000010111011010001110000000010;
				12'hC2B: data <= 32'b00000010111100000000101010010101;
				12'hC2C: data <= 32'b00000010111100101111110000011000;
				12'hC2D: data <= 32'b00000010111101011111000010001110;
				12'hC2E: data <= 32'b00000010111110001110011111111010;
				12'hC2F: data <= 32'b00000010111110111110001001011111;
				12'hC30: data <= 32'b00000010111111101101111111000000;
				12'hC31: data <= 32'b00000011000000011110000000100000;
				12'hC32: data <= 32'b00000011000001001110001110000001;
				12'hC33: data <= 32'b00000011000001111110100111101000;
				12'hC34: data <= 32'b00000011000010101111001101010110;
				12'hC35: data <= 32'b00000011000011011111111111010000;
				12'hC36: data <= 32'b00000011000100010000111101010111;
				12'hC37: data <= 32'b00000011000101000010000111101111;
				12'hC38: data <= 32'b00000011000101110011011110011100;
				12'hC39: data <= 32'b00000011000110100101000001100000;
				12'hC3A: data <= 32'b00000011000111010110110000111110;
				12'hC3B: data <= 32'b00000011001000001000101100111001;
				12'hC3C: data <= 32'b00000011001000111010110101010101;
				12'hC3D: data <= 32'b00000011001001101101001010010101;
				12'hC3E: data <= 32'b00000011001010011111101011111011;
				12'hC3F: data <= 32'b00000011001011010010011010001100;
				12'hC40: data <= 32'b00000011001100000101010101001001;
				12'hC41: data <= 32'b00000011001100111000011100110111;
				12'hC42: data <= 32'b00000011001101101011110001011001;
				12'hC43: data <= 32'b00000011001110011111010010110001;
				12'hC44: data <= 32'b00000011001111010011000001000011;
				12'hC45: data <= 32'b00000011010000000110111100010011;
				12'hC46: data <= 32'b00000011010000111011000100100011;
				12'hC47: data <= 32'b00000011010001101111011001110110;
				12'hC48: data <= 32'b00000011010010100011111100010001;
				12'hC49: data <= 32'b00000011010011011000101011110101;
				12'hC4A: data <= 32'b00000011010100001101101000101000;
				12'hC4B: data <= 32'b00000011010101000010110010101011;
				12'hC4C: data <= 32'b00000011010101111000001010000010;
				12'hC4D: data <= 32'b00000011010110101101101110110001;
				12'hC4E: data <= 32'b00000011010111100011100000111011;
				12'hC4F: data <= 32'b00000011011000011001100000100011;
				12'hC50: data <= 32'b00000011011001001111101101101100;
				12'hC51: data <= 32'b00000011011010000110001000011011;
				12'hC52: data <= 32'b00000011011010111100110000110001;
				12'hC53: data <= 32'b00000011011011110011100110110100;
				12'hC54: data <= 32'b00000011011100101010101010100110;
				12'hC55: data <= 32'b00000011011101100001111100001011;
				12'hC56: data <= 32'b00000011011110011001011011100101;
				12'hC57: data <= 32'b00000011011111010001001000111001;
				12'hC58: data <= 32'b00000011100000001001000100001011;
				12'hC59: data <= 32'b00000011100001000001001101011101;
				12'hC5A: data <= 32'b00000011100001111001100100110011;
				12'hC5B: data <= 32'b00000011100010110010001010010000;
				12'hC5C: data <= 32'b00000011100011101010111101111001;
				12'hC5D: data <= 32'b00000011100100100011111111110000;
				12'hC5E: data <= 32'b00000011100101011101001111111010;
				12'hC5F: data <= 32'b00000011100110010110101110011010;
				12'hC60: data <= 32'b00000011100111010000011011010010;
				12'hC61: data <= 32'b00000011101000001010010110101000;
				12'hC62: data <= 32'b00000011101001000100100000011111;
				12'hC63: data <= 32'b00000011101001111110111000111010;
				12'hC64: data <= 32'b00000011101010111001011111111101;
				12'hC65: data <= 32'b00000011101011110100010101101011;
				12'hC66: data <= 32'b00000011101100101111011010001001;
				12'hC67: data <= 32'b00000011101101101010101101011001;
				12'hC68: data <= 32'b00000011101110100110001111100001;
				12'hC69: data <= 32'b00000011101111100010000000100010;
				12'hC6A: data <= 32'b00000011110000011110000000100010;
				12'hC6B: data <= 32'b00000011110001011010001111100100;
				12'hC6C: data <= 32'b00000011110010010110101101101011;
				12'hC6D: data <= 32'b00000011110011010011011010111100;
				12'hC6E: data <= 32'b00000011110100010000010111011010;
				12'hC6F: data <= 32'b00000011110101001101100011001001;
				12'hC70: data <= 32'b00000011110110001010111110001101;
				12'hC71: data <= 32'b00000011110111001000101000101001;
				12'hC72: data <= 32'b00000011111000000110100010100010;
				12'hC73: data <= 32'b00000011111001000100101011111100;
				12'hC74: data <= 32'b00000011111010000011000100111010;
				12'hC75: data <= 32'b00000011111011000001101101100000;
				12'hC76: data <= 32'b00000011111100000000100101110010;
				12'hC77: data <= 32'b00000011111100111111101101110100;
				12'hC78: data <= 32'b00000011111101111111000101101010;
				12'hC79: data <= 32'b00000011111110111110101101011000;
				12'hC7A: data <= 32'b00000011111111111110100101000010;
				12'hC7B: data <= 32'b00000100000000111110101100101100;
				12'hC7C: data <= 32'b00000100000001111111000100011010;
				12'hC7D: data <= 32'b00000100000010111111101100001111;
				12'hC7E: data <= 32'b00000100000100000000100100010001;
				12'hC7F: data <= 32'b00000100000101000001101100100011;
				12'hC80: data <= 32'b00000100000110000011000101001001;
				12'hC81: data <= 32'b00000100000111000100101110000111;
				12'hC82: data <= 32'b00000100001000000110100111100001;
				12'hC83: data <= 32'b00000100001001001000110001011100;
				12'hC84: data <= 32'b00000100001010001011001011111011;
				12'hC85: data <= 32'b00000100001011001101110111000011;
				12'hC86: data <= 32'b00000100001100010000110010111000;
				12'hC87: data <= 32'b00000100001101010011111111011110;
				12'hC88: data <= 32'b00000100001110010111011100111001;
				12'hC89: data <= 32'b00000100001111011011001011001110;
				12'hC8A: data <= 32'b00000100010000011111001010100000;
				12'hC8B: data <= 32'b00000100010001100011011010110101;
				12'hC8C: data <= 32'b00000100010010100111111100001111;
				12'hC8D: data <= 32'b00000100010011101100101110110100;
				12'hC8E: data <= 32'b00000100010100110001110010101000;
				12'hC8F: data <= 32'b00000100010101110111000111101111;
				12'hC90: data <= 32'b00000100010110111100101110001101;
				12'hC91: data <= 32'b00000100011000000010100110001000;
				12'hC92: data <= 32'b00000100011001001000101111100010;
				12'hC93: data <= 32'b00000100011010001111001010100001;
				12'hC94: data <= 32'b00000100011011010101110111001001;
				12'hC95: data <= 32'b00000100011100011100110101011110;
				12'hC96: data <= 32'b00000100011101100100000101100101;
				12'hC97: data <= 32'b00000100011110101011100111100010;
				12'hC98: data <= 32'b00000100011111110011011011011010;
				12'hC99: data <= 32'b00000100100000111011100001010001;
				12'hC9A: data <= 32'b00000100100010000011111001001100;
				12'hC9B: data <= 32'b00000100100011001100100011010000;
				12'hC9C: data <= 32'b00000100100100010101011111100000;
				12'hC9D: data <= 32'b00000100100101011110101110000001;
				12'hC9E: data <= 32'b00000100100110101000001110111000;
				12'hC9F: data <= 32'b00000100100111110010000010001010;
				12'hCA0: data <= 32'b00000100101000111100000111111011;
				12'hCA1: data <= 32'b00000100101010000110100000001111;
				12'hCA2: data <= 32'b00000100101011010001001011001100;
				12'hCA3: data <= 32'b00000100101100011100001000110110;
				12'hCA4: data <= 32'b00000100101101100111011001010010;
				12'hCA5: data <= 32'b00000100101110110010111100100101;
				12'hCA6: data <= 32'b00000100101111111110110010110010;
				12'hCA7: data <= 32'b00000100110001001010111100000000;
				12'hCA8: data <= 32'b00000100110010010111011000010010;
				12'hCA9: data <= 32'b00000100110011100100000111101101;
				12'hCAA: data <= 32'b00000100110100110001001010010111;
				12'hCAB: data <= 32'b00000100110101111110100000010100;
				12'hCAC: data <= 32'b00000100110111001100001001101001;
				12'hCAD: data <= 32'b00000100111000011010000110011011;
				12'hCAE: data <= 32'b00000100111001101000010110101110;
				12'hCAF: data <= 32'b00000100111010110110111010101000;
				12'hCB0: data <= 32'b00000100111100000101110010001101;
				12'hCB1: data <= 32'b00000100111101010100111101100010;
				12'hCB2: data <= 32'b00000100111110100100011100101101;
				12'hCB3: data <= 32'b00000100111111110100001111110010;
				12'hCB4: data <= 32'b00000101000001000100010110110111;
				12'hCB5: data <= 32'b00000101000010010100110010000000;
				12'hCB6: data <= 32'b00000101000011100101100001010001;
				12'hCB7: data <= 32'b00000101000100110110100100110010;
				12'hCB8: data <= 32'b00000101000110000111111100100110;
				12'hCB9: data <= 32'b00000101000111011001101000110010;
				12'hCBA: data <= 32'b00000101001000101011101001011100;
				12'hCBB: data <= 32'b00000101001001111101111110101000;
				12'hCBC: data <= 32'b00000101001011010000101000011101;
				12'hCBD: data <= 32'b00000101001100100011100110111110;
				12'hCBE: data <= 32'b00000101001101110110111010010010;
				12'hCBF: data <= 32'b00000101001111001010100010011101;
				12'hCC0: data <= 32'b00000101010000011110011111100101;
				12'hCC1: data <= 32'b00000101010001110010110001101111;
				12'hCC2: data <= 32'b00000101010011000111011001000000;
				12'hCC3: data <= 32'b00000101010100011100010101011101;
				12'hCC4: data <= 32'b00000101010101110001100111001100;
				12'hCC5: data <= 32'b00000101010111000111001110010010;
				12'hCC6: data <= 32'b00000101011000011101001010110101;
				12'hCC7: data <= 32'b00000101011001110011011100111001;
				12'hCC8: data <= 32'b00000101011011001010000100100101;
				12'hCC9: data <= 32'b00000101011100100001000001111110;
				12'hCCA: data <= 32'b00000101011101111000010101001000;
				12'hCCB: data <= 32'b00000101011111001111111110001010;
				12'hCCC: data <= 32'b00000101100000100111111101001001;
				12'hCCD: data <= 32'b00000101100010000000010010001010;
				12'hCCE: data <= 32'b00000101100011011000111101010100;
				12'hCCF: data <= 32'b00000101100100110001111110101011;
				12'hCD0: data <= 32'b00000101100110001011010110010101;
				12'hCD1: data <= 32'b00000101100111100101000100011000;
				12'hCD2: data <= 32'b00000101101000111111001000111001;
				12'hCD3: data <= 32'b00000101101010011001100011111110;
				12'hCD4: data <= 32'b00000101101011110100010101101101;
				12'hCD5: data <= 32'b00000101101101001111011110001011;
				12'hCD6: data <= 32'b00000101101110101010111101011110;
				12'hCD7: data <= 32'b00000101110000000110110011101100;
				12'hCD8: data <= 32'b00000101110001100011000000111010;
				12'hCD9: data <= 32'b00000101110010111111100101001110;
				12'hCDA: data <= 32'b00000101110100011100100000101110;
				12'hCDB: data <= 32'b00000101110101111001110011100000;
				12'hCDC: data <= 32'b00000101110111010111011101101010;
				12'hCDD: data <= 32'b00000101111000110101011111010001;
				12'hCDE: data <= 32'b00000101111010010011111000011100;
				12'hCDF: data <= 32'b00000101111011110010101001001111;
				12'hCE0: data <= 32'b00000101111101010001110001110010;
				12'hCE1: data <= 32'b00000101111110110001010010001010;
				12'hCE2: data <= 32'b00000110000000010001001010011101;
				12'hCE3: data <= 32'b00000110000001110001011010110001;
				12'hCE4: data <= 32'b00000110000011010010000011001101;
				12'hCE5: data <= 32'b00000110000100110011000011110101;
				12'hCE6: data <= 32'b00000110000110010100011100110001;
				12'hCE7: data <= 32'b00000110000111110110001110000101;
				12'hCE8: data <= 32'b00000110001001011000010111111010;
				12'hCE9: data <= 32'b00000110001010111010111010010011;
				12'hCEA: data <= 32'b00000110001100011101110101011001;
				12'hCEB: data <= 32'b00000110001110000001001001010000;
				12'hCEC: data <= 32'b00000110001111100100110110000000;
				12'hCED: data <= 32'b00000110010001001000111011101101;
				12'hCEE: data <= 32'b00000110010010101101011010100000;
				12'hCEF: data <= 32'b00000110010100010010010010011101;
				12'hCF0: data <= 32'b00000110010101110111100011101011;
				12'hCF1: data <= 32'b00000110010111011101001110010001;
				12'hCF2: data <= 32'b00000110011001000011010010010100;
				12'hCF3: data <= 32'b00000110011010101001101111111100;
				12'hCF4: data <= 32'b00000110011100010000100111001110;
				12'hCF5: data <= 32'b00000110011101110111111000010010;
				12'hCF6: data <= 32'b00000110011111011111100011001101;
				12'hCF7: data <= 32'b00000110100001000111101000000101;
				12'hCF8: data <= 32'b00000110100010110000000111000011;
				12'hCF9: data <= 32'b00000110100100011001000000001011;
				12'hCFA: data <= 32'b00000110100110000010010011100101;
				12'hCFB: data <= 32'b00000110100111101100000001010111;
				12'hCFC: data <= 32'b00000110101001010110001001101000;
				12'hCFD: data <= 32'b00000110101011000000101100011110;
				12'hCFE: data <= 32'b00000110101100101011101010000000;
				12'hCFF: data <= 32'b00000110101110010111000010010101;
				12'hD00: data <= 32'b00000110110000000010110101100100;
				12'hD01: data <= 32'b00000110110001101111000011110010;
				12'hD02: data <= 32'b00000110110011011011101101001000;
				12'hD03: data <= 32'b00000110110101001000110001101011;
				12'hD04: data <= 32'b00000110110110110110010001100011;
				12'hD05: data <= 32'b00000110111000100100001100110110;
				12'hD06: data <= 32'b00000110111010010010100011101100;
				12'hD07: data <= 32'b00000110111100000001010110001011;
				12'hD08: data <= 32'b00000110111101110000100100011001;
				12'hD09: data <= 32'b00000110111111100000001110011111;
				12'hD0A: data <= 32'b00000111000001010000010100100011;
				12'hD0B: data <= 32'b00000111000011000000110110101100;
				12'hD0C: data <= 32'b00000111000100110001110101000001;
				12'hD0D: data <= 32'b00000111000110100011001111101001;
				12'hD0E: data <= 32'b00000111001000010101000110101011;
				12'hD0F: data <= 32'b00000111001010000111011010001110;
				12'hD10: data <= 32'b00000111001011111010001010011010;
				12'hD11: data <= 32'b00000111001101101101010111010110;
				12'hD12: data <= 32'b00000111001111100001000001001000;
				12'hD13: data <= 32'b00000111010001010101000111111001;
				12'hD14: data <= 32'b00000111010011001001101011101111;
				12'hD15: data <= 32'b00000111010100111110101100110001;
				12'hD16: data <= 32'b00000111010110110100001011000111;
				12'hD17: data <= 32'b00000111011000101010000110111001;
				12'hD18: data <= 32'b00000111011010100000100000001101;
				12'hD19: data <= 32'b00000111011100010111010111001100;
				12'hD1A: data <= 32'b00000111011110001110101011111011;
				12'hD1B: data <= 32'b00000111100000000110011110100100;
				12'hD1C: data <= 32'b00000111100001111110101111001101;
				12'hD1D: data <= 32'b00000111100011110111011101111110;
				12'hD1E: data <= 32'b00000111100101110000101010111111;
				12'hD1F: data <= 32'b00000111100111101010010110010110;
				12'hD20: data <= 32'b00000111101001100100100000001100;
				12'hD21: data <= 32'b00000111101011011111001000101001;
				12'hD22: data <= 32'b00000111101101011010001111110011;
				12'hD23: data <= 32'b00000111101111010101110101110011;
				12'hD24: data <= 32'b00000111110001010001111010110001;
				12'hD25: data <= 32'b00000111110011001110011110110011;
				12'hD26: data <= 32'b00000111110101001011100010000011;
				12'hD27: data <= 32'b00000111110111001001000100100111;
				12'hD28: data <= 32'b00000111111001000111000110101000;
				12'hD29: data <= 32'b00000111111011000101101000001101;
				12'hD2A: data <= 32'b00000111111101000100101001011111;
				12'hD2B: data <= 32'b00000111111111000100001010100100;
				12'hD2C: data <= 32'b00001000000001000100001011100110;
				12'hD2D: data <= 32'b00001000000011000100101100101101;
				12'hD2E: data <= 32'b00001000000101000101101110000000;
				12'hD2F: data <= 32'b00001000000111000111001111100111;
				12'hD30: data <= 32'b00001000001001001001010001101010;
				12'hD31: data <= 32'b00001000001011001011110100010010;
				12'hD32: data <= 32'b00001000001101001110110111100111;
				12'hD33: data <= 32'b00001000001111010010011011110001;
				12'hD34: data <= 32'b00001000010001010110100000111000;
				12'hD35: data <= 32'b00001000010011011011000111000100;
				12'hD36: data <= 32'b00001000010101100000001110011110;
				12'hD37: data <= 32'b00001000010111100101110111001110;
				12'hD38: data <= 32'b00001000011001101100000001011100;
				12'hD39: data <= 32'b00001000011011110010101101010001;
				12'hD3A: data <= 32'b00001000011101111001111010110110;
				12'hD3B: data <= 32'b00001000100000000001101010010010;
				12'hD3C: data <= 32'b00001000100010001001111011101110;
				12'hD3D: data <= 32'b00001000100100010010101111010010;
				12'hD3E: data <= 32'b00001000100110011100000101001000;
				12'hD3F: data <= 32'b00001000101000100101111101011000;
				12'hD40: data <= 32'b00001000101010110000011000001010;
				12'hD41: data <= 32'b00001000101100111011010101100111;
				12'hD42: data <= 32'b00001000101111000110110101110111;
				12'hD43: data <= 32'b00001000110001010010111001000101;
				12'hD44: data <= 32'b00001000110011011111011111010111;
				12'hD45: data <= 32'b00001000110101101100101000110111;
				12'hD46: data <= 32'b00001000110111111010010101101110;
				12'hD47: data <= 32'b00001000111010001000100110000101;
				12'hD48: data <= 32'b00001000111100010111011010000100;
				12'hD49: data <= 32'b00001000111110100110110001110101;
				12'hD4A: data <= 32'b00001001000000110110101101100000;
				12'hD4B: data <= 32'b00001001000011000111001101001111;
				12'hD4C: data <= 32'b00001001000101011000010001001010;
				12'hD4D: data <= 32'b00001001000111101001111001011010;
				12'hD4E: data <= 32'b00001001001001111100000110001010;
				12'hD4F: data <= 32'b00001001001100001110110111100001;
				12'hD50: data <= 32'b00001001001110100010001101101000;
				12'hD51: data <= 32'b00001001010000110110001000101010;
				12'hD52: data <= 32'b00001001010011001010101000110000;
				12'hD53: data <= 32'b00001001010101011111101110000010;
				12'hD54: data <= 32'b00001001010111110101011000101010;
				12'hD55: data <= 32'b00001001011010001011101000110001;
				12'hD56: data <= 32'b00001001011100100010011110100010;
				12'hD57: data <= 32'b00001001011110111001111010000100;
				12'hD58: data <= 32'b00001001100001010001111011100010;
				12'hD59: data <= 32'b00001001100011101010100011000101;
				12'hD5A: data <= 32'b00001001100110000011110000110110;
				12'hD5B: data <= 32'b00001001101000011101100101000000;
				12'hD5C: data <= 32'b00001001101010110111111111101100;
				12'hD5D: data <= 32'b00001001101101010011000001000011;
				12'hD5E: data <= 32'b00001001101111101110101001010000;
				12'hD5F: data <= 32'b00001001110010001010111000011011;
				12'hD60: data <= 32'b00001001110100100111101110101111;
				12'hD61: data <= 32'b00001001110111000101001100010110;
				12'hD62: data <= 32'b00001001111001100011010001011001;
				12'hD63: data <= 32'b00001001111100000001111110000010;
				12'hD64: data <= 32'b00001001111110100001010010011011;
				12'hD65: data <= 32'b00001010000001000001001110101111;
				12'hD66: data <= 32'b00001010000011100001110011000110;
				12'hD67: data <= 32'b00001010000110000010111111101011;
				12'hD68: data <= 32'b00001010001000100100110100101001;
				12'hD69: data <= 32'b00001010001011000111010010001001;
				12'hD6A: data <= 32'b00001010001101101010011000010110;
				12'hD6B: data <= 32'b00001010010000001110000111011001;
				12'hD6C: data <= 32'b00001010010010110010011111011101;
				12'hD6D: data <= 32'b00001010010101010111100000101100;
				12'hD6E: data <= 32'b00001010010111111101001011010000;
				12'hD6F: data <= 32'b00001010011010100011011111010101;
				12'hD70: data <= 32'b00001010011101001010011101000100;
				12'hD71: data <= 32'b00001010011111110010000100100111;
				12'hD72: data <= 32'b00001010100010011010010110001001;
				12'hD73: data <= 32'b00001010100101000011010001110110;
				12'hD74: data <= 32'b00001010100111101100110111110110;
				12'hD75: data <= 32'b00001010101010010111001000010101;
				12'hD76: data <= 32'b00001010101101000010000011011110;
				12'hD77: data <= 32'b00001010101111101101101001011010;
				12'hD78: data <= 32'b00001010110010011001111010010110;
				12'hD79: data <= 32'b00001010110101000110110110011011;
				12'hD7A: data <= 32'b00001010110111110100011101110101;
				12'hD7B: data <= 32'b00001010111010100010110000101110;
				12'hD7C: data <= 32'b00001010111101010001101111010001;
				12'hD7D: data <= 32'b00001011000000000001011001101001;
				12'hD7E: data <= 32'b00001011000010110001110000000001;
				12'hD7F: data <= 32'b00001011000101100010110010100101;
				12'hD80: data <= 32'b00001011001000010100100001011110;
				12'hD81: data <= 32'b00001011001011000110111100111001;
				12'hD82: data <= 32'b00001011001101111010000101000000;
				12'hD83: data <= 32'b00001011010000101101111001111111;
				12'hD84: data <= 32'b00001011010011100010011100000001;
				12'hD85: data <= 32'b00001011010110010111101011010001;
				12'hD86: data <= 32'b00001011011001001101100111111011;
				12'hD87: data <= 32'b00001011011100000100010010001001;
				12'hD88: data <= 32'b00001011011110111011101010000111;
				12'hD89: data <= 32'b00001011100001110011110000000010;
				12'hD8A: data <= 32'b00001011100100101100100100000011;
				12'hD8B: data <= 32'b00001011100111100110000110011000;
				12'hD8C: data <= 32'b00001011101010100000010111001010;
				12'hD8D: data <= 32'b00001011101101011011010110100111;
				12'hD8E: data <= 32'b00001011110000010111000100111010;
				12'hD8F: data <= 32'b00001011110011010011100010001101;
				12'hD90: data <= 32'b00001011110110010000101110101111;
				12'hD91: data <= 32'b00001011111001001110101010101001;
				12'hD92: data <= 32'b00001011111100001101010110001000;
				12'hD93: data <= 32'b00001011111111001100110001011000;
				12'hD94: data <= 32'b00001100000010001100111100100101;
				12'hD95: data <= 32'b00001100000101001101110111111010;
				12'hD96: data <= 32'b00001100001000001111100011100101;
				12'hD97: data <= 32'b00001100001011010001111111110000;
				12'hD98: data <= 32'b00001100001110010101001100101000;
				12'hD99: data <= 32'b00001100010001011001001010011010;
				12'hD9A: data <= 32'b00001100010100011101111001010010;
				12'hD9B: data <= 32'b00001100010111100011011001011011;
				12'hD9C: data <= 32'b00001100011010101001101011000011;
				12'hD9D: data <= 32'b00001100011101110000101110010101;
				12'hD9E: data <= 32'b00001100100000111000100011011110;
				12'hD9F: data <= 32'b00001100100100000001001010101011;
				12'hDA0: data <= 32'b00001100100111001010100100000111;
				12'hDA1: data <= 32'b00001100101010010100110000000001;
				12'hDA2: data <= 32'b00001100101101011111101110100100;
				12'hDA3: data <= 32'b00001100110000101011011111111100;
				12'hDA4: data <= 32'b00001100110011111000000100011000;
				12'hDA5: data <= 32'b00001100110111000101011100000011;
				12'hDA6: data <= 32'b00001100111010010011100111001010;
				12'hDA7: data <= 32'b00001100111101100010100101111011;
				12'hDA8: data <= 32'b00001101000000110010011000100010;
				12'hDA9: data <= 32'b00001101000100000010111111001011;
				12'hDAA: data <= 32'b00001101000111010100011010000101;
				12'hDAB: data <= 32'b00001101001010100110101001011101;
				12'hDAC: data <= 32'b00001101001101111001101101011111;
				12'hDAD: data <= 32'b00001101010001001101100110011000;
				12'hDAE: data <= 32'b00001101010100100010010100010110;
				12'hDAF: data <= 32'b00001101010111110111110111100111;
				12'hDB0: data <= 32'b00001101011011001110010000010110;
				12'hDB1: data <= 32'b00001101011110100101011110110011;
				12'hDB2: data <= 32'b00001101100001111101100011001010;
				12'hDB3: data <= 32'b00001101100101010110011101101001;
				12'hDB4: data <= 32'b00001101101000110000001110011110;
				12'hDB5: data <= 32'b00001101101100001010110101110101;
				12'hDB6: data <= 32'b00001101101111100110010011111101;
				12'hDB7: data <= 32'b00001101110011000010101001000100;
				12'hDB8: data <= 32'b00001101110110011111110101010110;
				12'hDB9: data <= 32'b00001101111001111101111001000011;
				12'hDBA: data <= 32'b00001101111101011100110100011000;
				12'hDBB: data <= 32'b00001110000000111100100111100010;
				12'hDBC: data <= 32'b00001110000100011101010010110000;
				12'hDBD: data <= 32'b00001110000111111110110110010000;
				12'hDBE: data <= 32'b00001110001011100001010010010000;
				12'hDBF: data <= 32'b00001110001111000100100110111110;
				12'hDC0: data <= 32'b00001110010010101000110100101000;
				12'hDC1: data <= 32'b00001110010110001101111011011101;
				12'hDC2: data <= 32'b00001110011001110011111011101011;
				12'hDC3: data <= 32'b00001110011101011010110101011111;
				12'hDC4: data <= 32'b00001110100001000010101001001010;
				12'hDC5: data <= 32'b00001110100100101011010110111001;
				12'hDC6: data <= 32'b00001110101000010100111110111010;
				12'hDC7: data <= 32'b00001110101011111111100001011101;
				12'hDC8: data <= 32'b00001110101111101010111110110000;
				12'hDC9: data <= 32'b00001110110011010111010111000010;
				12'hDCA: data <= 32'b00001110110111000100101010100000;
				12'hDCB: data <= 32'b00001110111010110010111001011100;
				12'hDCC: data <= 32'b00001110111110100010000100000010;
				12'hDCD: data <= 32'b00001111000010010010001010100011;
				12'hDCE: data <= 32'b00001111000110000011001101001100;
				12'hDCF: data <= 32'b00001111001001110101001100001110;
				12'hDD0: data <= 32'b00001111001101101000000111111000;
				12'hDD1: data <= 32'b00001111010001011100000000010111;
				12'hDD2: data <= 32'b00001111010101010000110101111101;
				12'hDD3: data <= 32'b00001111011001000110101000110111;
				12'hDD4: data <= 32'b00001111011100111101011001010110;
				12'hDD5: data <= 32'b00001111100000110101000111101001;
				12'hDD6: data <= 32'b00001111100100101101110011111111;
				12'hDD7: data <= 32'b00001111101000100111011110101000;
				12'hDD8: data <= 32'b00001111101100100010000111110100;
				12'hDD9: data <= 32'b00001111110000011101101111110010;
				12'hDDA: data <= 32'b00001111110100011010010110110001;
				12'hDDB: data <= 32'b00001111111000010111111101000010;
				12'hDDC: data <= 32'b00001111111100010110100010110101;
				12'hDDD: data <= 32'b00010000000000010110001000011001;
				12'hDDE: data <= 32'b00010000000100010110101101111110;
				12'hDDF: data <= 32'b00010000001000011000010011110101;
				12'hDE0: data <= 32'b00010000001100011010111010001110;
				12'hDE1: data <= 32'b00010000010000011110100001011000;
				12'hDE2: data <= 32'b00010000010100100011001001100100;
				12'hDE3: data <= 32'b00010000011000101000110011000010;
				12'hDE4: data <= 32'b00010000011100101111011110000011;
				12'hDE5: data <= 32'b00010000100000110111001010110111;
				12'hDE6: data <= 32'b00010000100100111111111001101110;
				12'hDE7: data <= 32'b00010000101001001001101010111001;
				12'hDE8: data <= 32'b00010000101101010100011110101001;
				12'hDE9: data <= 32'b00010000110001100000010101001110;
				12'hDEA: data <= 32'b00010000110101101101001110111001;
				12'hDEB: data <= 32'b00010000111001111011001011111011;
				12'hDEC: data <= 32'b00010000111110001010001100100101;
				12'hDED: data <= 32'b00010001000010011010010001000111;
				12'hDEE: data <= 32'b00010001000110101011011001110011;
				12'hDEF: data <= 32'b00010001001010111101100110111010;
				12'hDF0: data <= 32'b00010001001111010000111000101100;
				12'hDF1: data <= 32'b00010001010011100101001111011100;
				12'hDF2: data <= 32'b00010001010111111010101011011010;
				12'hDF3: data <= 32'b00010001011100010001001100110111;
				12'hDF4: data <= 32'b00010001100000101000110100000110;
				12'hDF5: data <= 32'b00010001100101000001100001010111;
				12'hDF6: data <= 32'b00010001101001011011010100111100;
				12'hDF7: data <= 32'b00010001101101110110001111000111;
				12'hDF8: data <= 32'b00010001110010010010010000001010;
				12'hDF9: data <= 32'b00010001110110101111011000010101;
				12'hDFA: data <= 32'b00010001111011001101100111111100;
				12'hDFB: data <= 32'b00010001111111101100111111001111;
				12'hDFC: data <= 32'b00010010000100001101011110100010;
				12'hDFD: data <= 32'b00010010001000101111000110000101;
				12'hDFE: data <= 32'b00010010001101010001110110001011;
				12'hDFF: data <= 32'b00010010010001110101101111000110;
				12'hE00: data <= 32'b00010010010110011010110001001000;
				12'hE01: data <= 32'b00010010011011000000111100100100;
				12'hE02: data <= 32'b00010010011111101000010001101101;
				12'hE03: data <= 32'b00010010100100010000110000110011;
				12'hE04: data <= 32'b00010010101000111010011010001011;
				12'hE05: data <= 32'b00010010101101100101001110000111;
				12'hE06: data <= 32'b00010010110010010001001100111001;
				12'hE07: data <= 32'b00010010110110111110010110110011;
				12'hE08: data <= 32'b00010010111011101100101100001010;
				12'hE09: data <= 32'b00010011000000011100001101010000;
				12'hE0A: data <= 32'b00010011000101001100111010010111;
				12'hE0B: data <= 32'b00010011001001111110110011110011;
				12'hE0C: data <= 32'b00010011001110110001111001111000;
				12'hE0D: data <= 32'b00010011010011100110001100110111;
				12'hE0E: data <= 32'b00010011011000011011101101000100;
				12'hE0F: data <= 32'b00010011011101010010011010110100;
				12'hE10: data <= 32'b00010011100010001010010110011000;
				12'hE11: data <= 32'b00010011100111000011100000000101;
				12'hE12: data <= 32'b00010011101011111101111000001111;
				12'hE13: data <= 32'b00010011110000111001011111001000;
				12'hE14: data <= 32'b00010011110101110110010101000101;
				12'hE15: data <= 32'b00010011111010110100011010011001;
				12'hE16: data <= 32'b00010011111111110011101111011001;
				12'hE17: data <= 32'b00010100000100110100010100011000;
				12'hE18: data <= 32'b00010100001001110110001001101010;
				12'hE19: data <= 32'b00010100001110111001001111100011;
				12'hE1A: data <= 32'b00010100010011111101100110011000;
				12'hE1B: data <= 32'b00010100011001000011001110011101;
				12'hE1C: data <= 32'b00010100011110001010001000000110;
				12'hE1D: data <= 32'b00010100100011010010010011101000;
				12'hE1E: data <= 32'b00010100101000011011110001010111;
				12'hE1F: data <= 32'b00010100101101100110100001101000;
				12'hE20: data <= 32'b00010100110010110010100100101111;
				12'hE21: data <= 32'b00010100110111111111111011000001;
				12'hE22: data <= 32'b00010100111101001110100100110011;
				12'hE23: data <= 32'b00010101000010011110100010011010;
				12'hE24: data <= 32'b00010101000111101111110100001011;
				12'hE25: data <= 32'b00010101001101000010011010011011;
				12'hE26: data <= 32'b00010101010010010110010101100000;
				12'hE27: data <= 32'b00010101010111101011100101101101;
				12'hE28: data <= 32'b00010101011101000010001011011010;
				12'hE29: data <= 32'b00010101100010011010000110111010;
				12'hE2A: data <= 32'b00010101100111110011011000100100;
				12'hE2B: data <= 32'b00010101101101001110000000101110;
				12'hE2C: data <= 32'b00010101110010101001111111101100;
				12'hE2D: data <= 32'b00010101111000000111010101110101;
				12'hE2E: data <= 32'b00010101111101100110000011011110;
				12'hE2F: data <= 32'b00010110000011000110001000111110;
				12'hE30: data <= 32'b00010110001000100111100110101010;
				12'hE31: data <= 32'b00010110001110001010011100111001;
				12'hE32: data <= 32'b00010110010011101110101100000000;
				12'hE33: data <= 32'b00010110011001010100010100010110;
				12'hE34: data <= 32'b00010110011110111011010110010001;
				12'hE35: data <= 32'b00010110100100100011110010001001;
				12'hE36: data <= 32'b00010110101010001101101000010010;
				12'hE37: data <= 32'b00010110101111111000111001000100;
				12'hE38: data <= 32'b00010110110101100101100100110110;
				12'hE39: data <= 32'b00010110111011010011101011111110;
				12'hE3A: data <= 32'b00010111000001000011001110110100;
				12'hE3B: data <= 32'b00010111000110110100001101101101;
				12'hE3C: data <= 32'b00010111001100100110101001000010;
				12'hE3D: data <= 32'b00010111010010011010100001001010;
				12'hE3E: data <= 32'b00010111011000001111110110011011;
				12'hE3F: data <= 32'b00010111011110000110101001001101;
				12'hE40: data <= 32'b00010111100011111110111001110111;
				12'hE41: data <= 32'b00010111101001111000101000110001;
				12'hE42: data <= 32'b00010111101111110011110110010011;
				12'hE43: data <= 32'b00010111110101110000100010110101;
				12'hE44: data <= 32'b00010111111011101110101110101101;
				12'hE45: data <= 32'b00011000000001101110011010010100;
				12'hE46: data <= 32'b00011000000111101111100110000010;
				12'hE47: data <= 32'b00011000001101110010010010001111;
				12'hE48: data <= 32'b00011000010011110110011111010011;
				12'hE49: data <= 32'b00011000011001111100001101100111;
				12'hE4A: data <= 32'b00011000100000000011011101100010;
				12'hE4B: data <= 32'b00011000100110001100001111011110;
				12'hE4C: data <= 32'b00011000101100010110100011110010;
				12'hE4D: data <= 32'b00011000110010100010011010111000;
				12'hE4E: data <= 32'b00011000111000101111110101001000;
				12'hE4F: data <= 32'b00011000111110111110110010111011;
				12'hE50: data <= 32'b00011001000101001111010100101001;
				12'hE51: data <= 32'b00011001001011100001011010101101;
				12'hE52: data <= 32'b00011001010001110101000101011111;
				12'hE53: data <= 32'b00011001011000001010010101011000;
				12'hE54: data <= 32'b00011001011110100001001010110010;
				12'hE55: data <= 32'b00011001100100111001100110000110;
				12'hE56: data <= 32'b00011001101011010011100111101110;
				12'hE57: data <= 32'b00011001110001101111010000000011;
				12'hE58: data <= 32'b00011001111000001100011111011111;
				12'hE59: data <= 32'b00011001111110101011010110011011;
				12'hE5A: data <= 32'b00011010000101001011110101010010;
				12'hE5B: data <= 32'b00011010001011101101111100011110;
				12'hE5C: data <= 32'b00011010010010010001101100011001;
				12'hE5D: data <= 32'b00011010011000110111000101011101;
				12'hE5E: data <= 32'b00011010011111011110001000000101;
				12'hE5F: data <= 32'b00011010100110000110110100101010;
				12'hE60: data <= 32'b00011010101100110001001011101000;
				12'hE61: data <= 32'b00011010110011011101001101011001;
				12'hE62: data <= 32'b00011010111010001010111010011000;
				12'hE63: data <= 32'b00011011000000111010010010111111;
				12'hE64: data <= 32'b00011011000111101011010111101010;
				12'hE65: data <= 32'b00011011001110011110001000110100;
				12'hE66: data <= 32'b00011011010101010010100110111000;
				12'hE67: data <= 32'b00011011011100001000110010010001;
				12'hE68: data <= 32'b00011011100011000000101011011010;
				12'hE69: data <= 32'b00011011101001111010010010101111;
				12'hE6A: data <= 32'b00011011110000110101101000101101;
				12'hE6B: data <= 32'b00011011110111110010101101101101;
				12'hE6C: data <= 32'b00011011111110110001100010001101;
				12'hE6D: data <= 32'b00011100000101110010000110101000;
				12'hE6E: data <= 32'b00011100001100110100011011011001;
				12'hE6F: data <= 32'b00011100010011111000100000111111;
				12'hE70: data <= 32'b00011100011010111110010111110011;
				12'hE71: data <= 32'b00011100100010000110000000010100;
				12'hE72: data <= 32'b00011100101001001111011010111101;
				12'hE73: data <= 32'b00011100110000011010101000001011;
				12'hE74: data <= 32'b00011100110111100111101000011011;
				12'hE75: data <= 32'b00011100111110110110011100001001;
				12'hE76: data <= 32'b00011101000110000111000011110010;
				12'hE77: data <= 32'b00011101001101011001011111110100;
				12'hE78: data <= 32'b00011101010100101101110000101100;
				12'hE79: data <= 32'b00011101011100000011110110110111;
				12'hE7A: data <= 32'b00011101100011011011110010110001;
				12'hE7B: data <= 32'b00011101101010110101100100111010;
				12'hE7C: data <= 32'b00011101110010010001001101101110;
				12'hE7D: data <= 32'b00011101111001101110101101101011;
				12'hE7E: data <= 32'b00011110000001001110000101001110;
				12'hE7F: data <= 32'b00011110001000101111010100110111;
				12'hE80: data <= 32'b00011110010000010010011101000011;
				12'hE81: data <= 32'b00011110010111110111011110010000;
				12'hE82: data <= 32'b00011110011111011110011000111100;
				12'hE83: data <= 32'b00011110100111000111001101100110;
				12'hE84: data <= 32'b00011110101110110001111100101101;
				12'hE85: data <= 32'b00011110110110011110100110101111;
				12'hE86: data <= 32'b00011110111110001101001100001011;
				12'hE87: data <= 32'b00011111000101111101101101100000;
				12'hE88: data <= 32'b00011111001101110000001011001100;
				12'hE89: data <= 32'b00011111010101100100100101110000;
				12'hE8A: data <= 32'b00011111011101011010111101101001;
				12'hE8B: data <= 32'b00011111100101010011010011011001;
				12'hE8C: data <= 32'b00011111101101001101100111011110;
				12'hE8D: data <= 32'b00011111110101001001111010010111;
				12'hE8E: data <= 32'b00011111111101001000001100100101;
				12'hE8F: data <= 32'b00100000000101001000011110101000;
				12'hE90: data <= 32'b00100000001101001010110000111111;
				12'hE91: data <= 32'b00100000010101001111000100001011;
				12'hE92: data <= 32'b00100000011101010101011000101100;
				12'hE93: data <= 32'b00100000100101011101101111000010;
				12'hE94: data <= 32'b00100000101101101000000111101111;
				12'hE95: data <= 32'b00100000110101110100100011010001;
				12'hE96: data <= 32'b00100000111110000011000010001011;
				12'hE97: data <= 32'b00100001000110010011100100111101;
				12'hE98: data <= 32'b00100001001110100110001100001001;
				12'hE99: data <= 32'b00100001010110111010111000001110;
				12'hE9A: data <= 32'b00100001011111010001101001110000;
				12'hE9B: data <= 32'b00100001100111101010100001001111;
				12'hE9C: data <= 32'b00100001110000000101011111001100;
				12'hE9D: data <= 32'b00100001111000100010100100001001;
				12'hE9E: data <= 32'b00100010000001000001110000101001;
				12'hE9F: data <= 32'b00100010001001100011000101001101;
				12'hEA0: data <= 32'b00100010010010000110100010010111;
				12'hEA1: data <= 32'b00100010011010101100001000101010;
				12'hEA2: data <= 32'b00100010100011010011111000100111;
				12'hEA3: data <= 32'b00100010101011111101110010110001;
				12'hEA4: data <= 32'b00100010110100101001110111101100;
				12'hEA5: data <= 32'b00100010111101011000000111111001;
				12'hEA6: data <= 32'b00100011000110001000100011111011;
				12'hEA7: data <= 32'b00100011001110111011001100010111;
				12'hEA8: data <= 32'b00100011010111110000000001101101;
				12'hEA9: data <= 32'b00100011100000100111000100100011;
				12'hEAA: data <= 32'b00100011101001100000010101011100;
				12'hEAB: data <= 32'b00100011110010011011110100111010;
				12'hEAC: data <= 32'b00100011111011011001100011100010;
				12'hEAD: data <= 32'b00100100000100011001100001111000;
				12'hEAE: data <= 32'b00100100001101011011110000011111;
				12'hEAF: data <= 32'b00100100010110100000001111111100;
				12'hEB0: data <= 32'b00100100011111100111000000110011;
				12'hEB1: data <= 32'b00100100101000110000000011101000;
				12'hEB2: data <= 32'b00100100110001111011011001000001;
				12'hEB3: data <= 32'b00100100111011001001000001100001;
				12'hEB4: data <= 32'b00100101000100011000111101101110;
				12'hEB5: data <= 32'b00100101001101101011001110001100;
				12'hEB6: data <= 32'b00100101010110111111110011100010;
				12'hEB7: data <= 32'b00100101100000010110101110010011;
				12'hEB8: data <= 32'b00100101101001101111111111000101;
				12'hEB9: data <= 32'b00100101110011001011100110011111;
				12'hEBA: data <= 32'b00100101111100101001100101000101;
				12'hEBB: data <= 32'b00100110000110001001111011011110;
				12'hEBC: data <= 32'b00100110001111101100101010001111;
				12'hEBD: data <= 32'b00100110011001010001110010000000;
				12'hEBE: data <= 32'b00100110100010111001010011010101;
				12'hEBF: data <= 32'b00100110101100100011001110110110;
				12'hEC0: data <= 32'b00100110110110001111100101001010;
				12'hEC1: data <= 32'b00100110111111111110010110110110;
				12'hEC2: data <= 32'b00100111001001101111100100100010;
				12'hEC3: data <= 32'b00100111010011100011001110110101;
				12'hEC4: data <= 32'b00100111011101011001010110010111;
				12'hEC5: data <= 32'b00100111100111010001111011101110;
				12'hEC6: data <= 32'b00100111110001001100111111100010;
				12'hEC7: data <= 32'b00100111111011001010100010011011;
				12'hEC8: data <= 32'b00101000000101001010100101000000;
				12'hEC9: data <= 32'b00101000001111001101000111111010;
				12'hECA: data <= 32'b00101000011001010010001011110010;
				12'hECB: data <= 32'b00101000100011011001110001001110;
				12'hECC: data <= 32'b00101000101101100011111000111000;
				12'hECD: data <= 32'b00101000110111110000100011011000;
				12'hECE: data <= 32'b00101001000001111111110001010111;
				12'hECF: data <= 32'b00101001001100010001100011011110;
				12'hED0: data <= 32'b00101001010110100101111010010110;
				12'hED1: data <= 32'b00101001100000111100110110101001;
				12'hED2: data <= 32'b00101001101011010110011001000000;
				12'hED3: data <= 32'b00101001110101110010100010000100;
				12'hED4: data <= 32'b00101010000000010001010010011111;
				12'hED5: data <= 32'b00101010001010110010101010111011;
				12'hED6: data <= 32'b00101010010101010110101100000010;
				12'hED7: data <= 32'b00101010011111111101010110011111;
				12'hED8: data <= 32'b00101010101010100110101010111100;
				12'hED9: data <= 32'b00101010110101010010101010000011;
				12'hEDA: data <= 32'b00101011000000000001010100011111;
				12'hEDB: data <= 32'b00101011001010110010101010111011;
				12'hEDC: data <= 32'b00101011010101100110101110000011;
				12'hEDD: data <= 32'b00101011100000011101011110100001;
				12'hEDE: data <= 32'b00101011101011010110111101000000;
				12'hEDF: data <= 32'b00101011110110010011001010001110;
				12'hEE0: data <= 32'b00101100000001010010000110110100;
				12'hEE1: data <= 32'b00101100001100010011110011100000;
				12'hEE2: data <= 32'b00101100010111011000010000111101;
				12'hEE3: data <= 32'b00101100100010011111011111110111;
				12'hEE4: data <= 32'b00101100101101101001100000111011;
				12'hEE5: data <= 32'b00101100111000110110010100110110;
				12'hEE6: data <= 32'b00101101000100000101111100010101;
				12'hEE7: data <= 32'b00101101001111011000011000000100;
				12'hEE8: data <= 32'b00101101011010101101101000110000;
				12'hEE9: data <= 32'b00101101100110000101101111000111;
				12'hEEA: data <= 32'b00101101110001100000101011110111;
				12'hEEB: data <= 32'b00101101111100111110011111101100;
				12'hEEC: data <= 32'b00101110001000011111001011010110;
				12'hEED: data <= 32'b00101110010100000010101111100001;
				12'hEEE: data <= 32'b00101110011111101001001100111101;
				12'hEEF: data <= 32'b00101110101011010010100100010111;
				12'hEF0: data <= 32'b00101110110110111110110110011111;
				12'hEF1: data <= 32'b00101111000010101110000100000010;
				12'hEF2: data <= 32'b00101111001110100000001101110001;
				12'hEF3: data <= 32'b00101111011010010101010100011001;
				12'hEF4: data <= 32'b00101111100110001101011000101011;
				12'hEF5: data <= 32'b00101111110010001000011011010101;
				12'hEF6: data <= 32'b00101111111110000110011101001000;
				12'hEF7: data <= 32'b00110000001010000111011110110100;
				12'hEF8: data <= 32'b00110000010110001011100001001000;
				12'hEF9: data <= 32'b00110000100010010010100100110100;
				12'hEFA: data <= 32'b00110000101110011100101010101010;
				12'hEFB: data <= 32'b00110000111010101001110011011010;
				12'hEFC: data <= 32'b00110001000110111001111111110100;
				12'hEFD: data <= 32'b00110001010011001101010000101010;
				12'hEFE: data <= 32'b00110001011111100011100110101101;
				12'hEFF: data <= 32'b00110001101011111101000010101110;
				12'hF00: data <= 32'b00110001111000011001100101011111;
				12'hF01: data <= 32'b00110010000100111001001111110001;
				12'hF02: data <= 32'b00110010010001011100000010010111;
				12'hF03: data <= 32'b00110010011110000001111110000011;
				12'hF04: data <= 32'b00110010101010101011000011100111;
				12'hF05: data <= 32'b00110010110111010111010011110110;
				12'hF06: data <= 32'b00110011000100000110101111100010;
				12'hF07: data <= 32'b00110011010000111001010111011111;
				12'hF08: data <= 32'b00110011011101101111001100011111;
				12'hF09: data <= 32'b00110011101010101000001111010110;
				12'hF0A: data <= 32'b00110011110111100100100000111000;
				12'hF0B: data <= 32'b00110100000100100100000001111000;
				12'hF0C: data <= 32'b00110100010001100110110011001010;
				12'hF0D: data <= 32'b00110100011110101100110101100011;
				12'hF0E: data <= 32'b00110100101011110110001001110110;
				12'hF0F: data <= 32'b00110100111001000010110000111001;
				12'hF10: data <= 32'b00110101000110010010101011100001;
				12'hF11: data <= 32'b00110101010011100101111010100001;
				12'hF12: data <= 32'b00110101100000111100011110110000;
				12'hF13: data <= 32'b00110101101110010110011001000010;
				12'hF14: data <= 32'b00110101111011110011101010001110;
				12'hF15: data <= 32'b00110110001001010100010011001001;
				12'hF16: data <= 32'b00110110010110111000010100101010;
				12'hF17: data <= 32'b00110110100100011111101111100110;
				12'hF18: data <= 32'b00110110110010001010100100110100;
				12'hF19: data <= 32'b00110110111111111000110101001010;
				12'hF1A: data <= 32'b00110111001101101010100001100001;
				12'hF1B: data <= 32'b00110111011011011111101010101101;
				12'hF1C: data <= 32'b00110111101001011000010001101000;
				12'hF1D: data <= 32'b00110111110111010100010111001001;
				12'hF1E: data <= 32'b00111000000101010011111100000111;
				12'hF1F: data <= 32'b00111000010011010111000001011010;
				12'hF20: data <= 32'b00111000100001011101100111111010;
				12'hF21: data <= 32'b00111000101111100111110000100000;
				12'hF22: data <= 32'b00111000111101110101011100000101;
				12'hF23: data <= 32'b00111001001100000110101011100001;
				12'hF24: data <= 32'b00111001011010011011011111101110;
				12'hF25: data <= 32'b00111001101000110011111001100100;
				12'hF26: data <= 32'b00111001110111001111111001111110;
				12'hF27: data <= 32'b00111010000101101111100001110101;
				12'hF28: data <= 32'b00111010010100010010110010000010;
				12'hF29: data <= 32'b00111010100010111001101011100001;
				12'hF2A: data <= 32'b00111010110001100100001111001100;
				12'hF2B: data <= 32'b00111011000000010010011101111100;
				12'hF2C: data <= 32'b00111011001111000100011000101110;
				12'hF2D: data <= 32'b00111011011101111010000000011100;
				12'hF2E: data <= 32'b00111011101100110011010110000010;
				12'hF2F: data <= 32'b00111011111011110000011010011011;
				12'hF30: data <= 32'b00111100001010110001001110100011;
				12'hF31: data <= 32'b00111100011001110101110011010111;
				12'hF32: data <= 32'b00111100101000111110001001110001;
				12'hF33: data <= 32'b00111100111000001010010010110000;
				12'hF34: data <= 32'b00111101000111011010001111001111;
				12'hF35: data <= 32'b00111101010110101110000000001100;
				12'hF36: data <= 32'b00111101100110000101100110100100;
				12'hF37: data <= 32'b00111101110101100001000011010100;
				12'hF38: data <= 32'b00111110000101000000010111011010;
				12'hF39: data <= 32'b00111110010100100011100011110100;
				12'hF3A: data <= 32'b00111110100100001010101001100000;
				12'hF3B: data <= 32'b00111110110011110101101001011110;
				12'hF3C: data <= 32'b00111111000011100100100100101010;
				12'hF3D: data <= 32'b00111111010011010111011100000101;
				12'hF3E: data <= 32'b00111111100011001110010000101101;
				12'hF3F: data <= 32'b00111111110011001001000011100011;
				12'hF40: data <= 32'b01000000000011000111110101100100;
				12'hF41: data <= 32'b01000000010011001010100111110011;
				12'hF42: data <= 32'b01000000100011010001011011001110;
				12'hF43: data <= 32'b01000000110011011100010000110110;
				12'hF44: data <= 32'b01000001000011101011001001101100;
				12'hF45: data <= 32'b01000001010011111110000110110000;
				12'hF46: data <= 32'b01000001100100010101001001000101;
				12'hF47: data <= 32'b01000001110100110000010001101011;
				12'hF48: data <= 32'b01000010000101001111100001100100;
				12'hF49: data <= 32'b01000010010101110010111001110010;
				12'hF4A: data <= 32'b01000010100110011010011011010111;
				12'hF4B: data <= 32'b01000010110111000110000111010101;
				12'hF4C: data <= 32'b01000011000111110101111110110001;
				12'hF4D: data <= 32'b01000011011000101010000010101011;
				12'hF4E: data <= 32'b01000011101001100010010100001000;
				12'hF4F: data <= 32'b01000011111010011110110100001100;
				12'hF50: data <= 32'b01000100001011011111100011111001;
				12'hF51: data <= 32'b01000100011100100100100100010100;
				12'hF52: data <= 32'b01000100101101101101110110100010;
				12'hF53: data <= 32'b01000100111110111011011011100111;
				12'hF54: data <= 32'b01000101010000001101010100100111;
				12'hF55: data <= 32'b01000101100001100011100010101000;
				12'hF56: data <= 32'b01000101110010111110000110101111;
				12'hF57: data <= 32'b01000110000100011101000010000011;
				12'hF58: data <= 32'b01000110010110000000010101101000;
				12'hF59: data <= 32'b01000110100111101000000010100101;
				12'hF5A: data <= 32'b01000110111001010100001010000001;
				12'hF5B: data <= 32'b01000111001011000100101101000010;
				12'hF5C: data <= 32'b01000111011100111001101100101111;
				12'hF5D: data <= 32'b01000111101110110011001010010000;
				12'hF5E: data <= 32'b01001000000000110001000110101100;
				12'hF5F: data <= 32'b01001000010010110011100011001011;
				12'hF60: data <= 32'b01001000100100111010100000110110;
				12'hF61: data <= 32'b01001000110111000110000000110100;
				12'hF62: data <= 32'b01001001001001010110000100001110;
				12'hF63: data <= 32'b01001001011011101010101100001110;
				12'hF64: data <= 32'b01001001101110000011111001111101;
				12'hF65: data <= 32'b01001010000000100001101110100100;
				12'hF66: data <= 32'b01001010010011000100001011001101;
				12'hF67: data <= 32'b01001010100101101011010001000010;
				12'hF68: data <= 32'b01001010111000010111000001001110;
				12'hF69: data <= 32'b01001011001011000111011100111100;
				12'hF6A: data <= 32'b01001011011101111100100101010110;
				12'hF6B: data <= 32'b01001011110000110110011011101000;
				12'hF6C: data <= 32'b01001100000011110101000000111101;
				12'hF6D: data <= 32'b01001100010110111000010110100001;
				12'hF6E: data <= 32'b01001100101010000000011101100001;
				12'hF6F: data <= 32'b01001100111101001101010111001010;
				12'hF70: data <= 32'b01001101010000011111000100100111;
				12'hF71: data <= 32'b01001101100011110101100111000110;
				12'hF72: data <= 32'b01001101110111010000111111110100;
				12'hF73: data <= 32'b01001110001010110001010000000000;
				12'hF74: data <= 32'b01001110011110010110011000110110;
				12'hF75: data <= 32'b01001110110010000000011011100110;
				12'hF76: data <= 32'b01001111000101101111011001011110;
				12'hF77: data <= 32'b01001111011001100011010011101101;
				12'hF78: data <= 32'b01001111101101011100001011100011;
				12'hF79: data <= 32'b01010000000001011010000010001110;
				12'hF7A: data <= 32'b01010000010101011100111000111110;
				12'hF7B: data <= 32'b01010000101001100100110001000101;
				12'hF7C: data <= 32'b01010000111101110001101011110010;
				12'hF7D: data <= 32'b01010001010010000011101010010110;
				12'hF7E: data <= 32'b01010001100110011010101110000010;
				12'hF7F: data <= 32'b01010001111010110110111000001000;
				12'hF80: data <= 32'b01010010001111011000001001111001;
				12'hF81: data <= 32'b01010010100011111110100100101000;
				12'hF82: data <= 32'b01010010111000101010001001100111;
				12'hF83: data <= 32'b01010011001101011010111010001001;
				12'hF84: data <= 32'b01010011100010010000110111100000;
				12'hF85: data <= 32'b01010011110111001100000011000000;
				12'hF86: data <= 32'b01010100001100001100011101111110;
				12'hF87: data <= 32'b01010100100001010010001001101011;
				12'hF88: data <= 32'b01010100110110011101000111011111;
				12'hF89: data <= 32'b01010101001011101101011000101011;
				12'hF8A: data <= 32'b01010101100001000010111110100111;
				12'hF8B: data <= 32'b01010101110110011101111010100111;
				12'hF8C: data <= 32'b01010110001011111110001110000001;
				12'hF8D: data <= 32'b01010110100001100011111010001011;
				12'hF8E: data <= 32'b01010110110111001111000000011011;
				12'hF8F: data <= 32'b01010111001100111111100010001000;
				12'hF90: data <= 32'b01010111100010110101100000101001;
				12'hF91: data <= 32'b01010111111000110000111101010110;
				12'hF92: data <= 32'b01011000001110110001111001100101;
				12'hF93: data <= 32'b01011000100100111000010110110000;
				12'hF94: data <= 32'b01011000111011000100010110001110;
				12'hF95: data <= 32'b01011001010001010101111001011001;
				12'hF96: data <= 32'b01011001100111101101000001101001;
				12'hF97: data <= 32'b01011001111110001001110000010111;
				12'hF98: data <= 32'b01011010010100101100000110111111;
				12'hF99: data <= 32'b01011010101011010100000110111001;
				12'hF9A: data <= 32'b01011011000010000001110001100000;
				12'hF9B: data <= 32'b01011011011000110101001000010000;
				12'hF9C: data <= 32'b01011011101111101110001100100011;
				12'hF9D: data <= 32'b01011100000110101100111111110101;
				12'hF9E: data <= 32'b01011100011101110001100011100010;
				12'hF9F: data <= 32'b01011100110100111011111001000110;
				12'hFA0: data <= 32'b01011101001100001100000001111101;
				12'hFA1: data <= 32'b01011101100011100001111111100110;
				12'hFA2: data <= 32'b01011101111010111101110011011100;
				12'hFA3: data <= 32'b01011110010010011111011110111111;
				12'hFA4: data <= 32'b01011110101010000111000011101011;
				12'hFA5: data <= 32'b01011111000001110100100011000000;
				12'hFA6: data <= 32'b01011111011001100111111110011100;
				12'hFA7: data <= 32'b01011111110001100001010111011111;
				12'hFA8: data <= 32'b01100000001001100000101111101000;
				12'hFA9: data <= 32'b01100000100001100110001000010111;
				12'hFAA: data <= 32'b01100000111001110001100011001100;
				12'hFAB: data <= 32'b01100001010010000011000001101001;
				12'hFAC: data <= 32'b01100001101010011010100101001110;
				12'hFAD: data <= 32'b01100010000010111000001111011100;
				12'hFAE: data <= 32'b01100010011011011100000001110110;
				12'hFAF: data <= 32'b01100010110100000101111101111110;
				12'hFB0: data <= 32'b01100011001100110110000101010110;
				12'hFB1: data <= 32'b01100011100101101100011001100001;
				12'hFB2: data <= 32'b01100011111110101000111100000100;
				12'hFB3: data <= 32'b01100100010111101011101110100001;
				12'hFB4: data <= 32'b01100100110000110100110010011101;
				12'hFB5: data <= 32'b01100101001010000100001001011100;
				12'hFB6: data <= 32'b01100101100011011001110101000011;
				12'hFB7: data <= 32'b01100101111100110101110110111000;
				12'hFB8: data <= 32'b01100110010110011000010000100000;
				12'hFB9: data <= 32'b01100110110000000001000011100010;
				12'hFBA: data <= 32'b01100111001001110000010001100100;
				12'hFBB: data <= 32'b01100111100011100101111100001110;
				12'hFBC: data <= 32'b01100111111101100010000101000101;
				12'hFBD: data <= 32'b01101000010111100100101101110011;
				12'hFBE: data <= 32'b01101000110001101101110111111111;
				12'hFBF: data <= 32'b01101001001011111101100101010010;
				12'hFC0: data <= 32'b01101001100110010011110111010100;
				12'hFC1: data <= 32'b01101010000000110000101111110001;
				12'hFC2: data <= 32'b01101010011011010100010000010000;
				12'hFC3: data <= 32'b01101010110101111110011010011100;
				12'hFC4: data <= 32'b01101011010000101111010000000001;
				12'hFC5: data <= 32'b01101011101011100110110010101000;
				12'hFC6: data <= 32'b01101100000110100101000011111110;
				12'hFC7: data <= 32'b01101100100001101010000101101110;
				12'hFC8: data <= 32'b01101100111100110101111001100101;
				12'hFC9: data <= 32'b01101101011000001000100001001111;
				12'hFCA: data <= 32'b01101101110011100001111110011010;
				12'hFCB: data <= 32'b01101110001111000010010010110011;
				12'hFCC: data <= 32'b01101110101010101001100000001000;
				12'hFCD: data <= 32'b01101111000110010111101000001000;
				12'hFCE: data <= 32'b01101111100010001100101100100001;
				12'hFCF: data <= 32'b01101111111110001000101111000011;
				12'hFD0: data <= 32'b01110000011010001011110001011110;
				12'hFD1: data <= 32'b01110000110110010101110101100001;
				12'hFD2: data <= 32'b01110001010010100110111100111110;
				12'hFD3: data <= 32'b01110001101110111111001001100110;
				12'hFD4: data <= 32'b01110010001011011110011101001001;
				12'hFD5: data <= 32'b01110010101000000100111001011010;
				12'hFD6: data <= 32'b01110011000100110010100000001100;
				12'hFD7: data <= 32'b01110011100001100111010011010001;
				12'hFD8: data <= 32'b01110011111110100011010100011100;
				12'hFD9: data <= 32'b01110100011011100110100101100010;
				12'hFDA: data <= 32'b01110100111000110001001000010110;
				12'hFDB: data <= 32'b01110101010110000010111110101101;
				12'hFDC: data <= 32'b01110101110011011100001010011100;
				12'hFDD: data <= 32'b01110110010000111100101101011001;
				12'hFDE: data <= 32'b01110110101110100100101001011010;
				12'hFDF: data <= 32'b01110111001100010100000000010110;
				12'hFE0: data <= 32'b01110111101010001010110100000010;
				12'hFE1: data <= 32'b01111000001000001001000110010111;
				12'hFE2: data <= 32'b01111000100110001110111001001101;
				12'hFE3: data <= 32'b01111001000100011100001110011100;
				12'hFE4: data <= 32'b01111001100010110001000111111101;
				12'hFE5: data <= 32'b01111010000001001101100111101001;
				12'hFE6: data <= 32'b01111010011111110001101111011001;
				12'hFE7: data <= 32'b01111010111110011101100001001001;
				12'hFE8: data <= 32'b01111011011101010000111110110011;
				12'hFE9: data <= 32'b01111011111100001100001010010010;
				12'hFEA: data <= 32'b01111100011011001111000101100001;
				12'hFEB: data <= 32'b01111100111010011001110010011110;
				12'hFEC: data <= 32'b01111101011001101100010011000100;
				12'hFED: data <= 32'b01111101111001000110101001010001;
				12'hFEE: data <= 32'b01111110011000101000110111000011;
				12'hFEF: data <= 32'b01111110111000010010111110010111;
				12'hFF0: data <= 32'b01111111011000000101000001001100;
				12'hFF1: data <= 32'b01111111110111111111000001100010;
				12'hFF2: data <= 32'b10000000011000000001000001011000;
				12'hFF3: data <= 32'b10000000111000001011000010101110;
				12'hFF4: data <= 32'b10000001011000011101000111100100;
				12'hFF5: data <= 32'b10000001111000110111010001111101;
				12'hFF6: data <= 32'b10000010011001011001100011111000;
				12'hFF7: data <= 32'b10000010111010000011111111011010;
				12'hFF8: data <= 32'b10000011011010110110100110100100;
				12'hFF9: data <= 32'b10000011111011110001011011011001;
				12'hFFA: data <= 32'b10000100011100110100011111111101;
				12'hFFB: data <= 32'b10000100111101111111110110010101;
				12'hFFC: data <= 32'b10000101011111010011100000100101;
				12'hFFD: data <= 32'b10000110000000101111100000110010;
				12'hFFE: data <= 32'b10000110100010010011111001000010;
				12'hFFF: data <= 32'b10000111000100000000101011011011;
			endcase
		end
	end

endmodule
