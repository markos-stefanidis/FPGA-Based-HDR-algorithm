module g_red_lut(
	input clk,
	input clk_en,
	input [4:0] pixel,
	
	output reg [11:0] data
);

	always@(posedge clk) begin
		if(clk_en) begin
			case(pixel)
				5'h00: data <= 12'b000000000000;
				5'h01: data <= 12'b000001110101;
				5'h02: data <= 12'b000011110110;
				5'h03: data <= 12'b000101111100;
				5'h04: data <= 12'b000111100011;
				5'h05: data <= 12'b001000101110;
				5'h06: data <= 12'b001001101100;
				5'h07: data <= 12'b001010100000;
				5'h08: data <= 12'b001011001100;
				5'h09: data <= 12'b001011110011;
				5'h0A: data <= 12'b001100010101;
				5'h0B: data <= 12'b001100110101;
				5'h0C: data <= 12'b001101010011;
				5'h0D: data <= 12'b001101110001;
				5'h0E: data <= 12'b001110001111;
				5'h0F: data <= 12'b001110101111;
				5'h10: data <= 12'b001111010000;
				5'h11: data <= 12'b001111110010;
				5'h12: data <= 12'b010000010100;
				5'h13: data <= 12'b010000110100;
				5'h14: data <= 12'b010001010011;
				5'h15: data <= 12'b010001101111;
				5'h16: data <= 12'b010010001001;
				5'h17: data <= 12'b010010100010;
				5'h18: data <= 12'b010010111010;
				5'h19: data <= 12'b010011010000;
				5'h1A: data <= 12'b010011100101;
				5'h1B: data <= 12'b010011111000;
				5'h1C: data <= 12'b010100001010;
				5'h1D: data <= 12'b010100011110;
				5'h1E: data <= 12'b010100110011;
				5'h1F: data <= 12'b010101001011;
			endcase
		end
	end

endmodule
